-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 10 2025 16:58:16

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    xor_out_stat : out std_logic;
    mosi_output : out std_logic;
    miso_input : in std_logic;
    xor_out_dyn : out std_logic;
    sel_output : out std_logic;
    s14 : out std_logic;
    s12 : out std_logic;
    clk_output : out std_logic;
    CLK : in std_logic;
    s13 : out std_logic;
    RST_N : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__12279\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \DYNCNF_i_0\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_49\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_38\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_34\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_35\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_36\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_37\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uCZ0\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_6c_0_0\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_6b_0_0\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_2_0_0\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_5_0_0\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_6_0_0\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_6dZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_6eZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_6fZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_3_0_0\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_4_0_0\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_16\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_17\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_33\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_48\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_30\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_71\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_31\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_32\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_72\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_41\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_39\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_40\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_12\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_13\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_3\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_2\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_11\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_14\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_4\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_5\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_6\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_7\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_8\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_9\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_10\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_1\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_6iZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_6jZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_6gZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_6hZ0Z_0\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_stat_cry_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_stat_cry_1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_stat_cry_2\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_stat_cry_3\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_stat_cry_4\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_stat_cry_5\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_15\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_14\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_22\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_20\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_21\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_18\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_19\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_25\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_26\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_29\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_23\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_24\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_27\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_28\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_47\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_73\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_74\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_75\ : std_logic;
signal \FSM_TEST_inst_slow.N_134_1_cascade_\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_15\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_87\ : std_logic;
signal \FSM_TEST_inst_slow.G_31_1\ : std_logic;
signal \FSM_TEST_inst_slow.counter_statlde_0_cascade_\ : std_logic;
signal \FSM_TEST_inst_slow.current_state_RNIR2L81Z0Z_1\ : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idle_cry_0\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idle_cry_1\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idle_cry_2\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idle_cry_3\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idle_cry_4\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idle_cry_5\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idle_cry_6\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idle_RNIHR3A2Z0Z_7\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idleZ0Z_1\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idleZ0Z_2\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idleZ0Z_5\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idleZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_slow.N_109_0\ : std_logic;
signal \FSM_TEST_inst_slow.counter_dinZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_slow.counter_dinZ1Z_1\ : std_logic;
signal \FSM_TEST_inst_slow.N_134_1_i\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idleZ0Z_4\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idleZ0Z_3\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_stat_cry_3_THRU_CO\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_stat_cry_4_THRU_CO\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_stat_cry_2_THRU_CO\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_statlde_0_cascade_\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2Z0Z_1_cascade_\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_statZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_stat_cry_0_THRU_CO\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2Z0Z_1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_stat_cry_1_THRU_CO\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_statZ0Z_2\ : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idle_cry_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idle_cry_1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idle_cry_2\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idle_cry_3\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idle_cry_4\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_13\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_81\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_46\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_4\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_1\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_2\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_3\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_80\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_42\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_70\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_45\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_76\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_77\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_43\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_44\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_78\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_79\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \FSM_TEST_inst_slow.counter_stat_cry_0\ : std_logic;
signal \FSM_TEST_inst_slow.counter_stat_cry_1\ : std_logic;
signal \FSM_TEST_inst_slow.counter_stat_cry_2\ : std_logic;
signal \FSM_TEST_inst_slow.counter_stat_cry_3\ : std_logic;
signal \FSM_TEST_inst_slow.counter_stat_cry_4\ : std_logic;
signal \FSM_TEST_inst_slow.counter_stat_cry_5\ : std_logic;
signal \FSM_TEST_inst_slow.counter_statZ0Z_6\ : std_logic;
signal \FSM_TEST_inst_slow.current_state_ns_0_a3_1_4_0_cascade_\ : std_logic;
signal \FSM_TEST_inst_slow.current_state_ns_0_a3_1_5_0\ : std_logic;
signal \FSM_TEST_inst_slow.counter_statZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_slow.counter_stat_cry_1_THRU_CO\ : std_logic;
signal \FSM_TEST_inst_slow.counter_statZ0Z_2\ : std_logic;
signal \FSM_TEST_inst_slow.counter_stat_cry_2_THRU_CO\ : std_logic;
signal \FSM_TEST_inst_slow.counter_statZ0Z_3\ : std_logic;
signal \FSM_TEST_inst_slow.counter_stat_cry_0_THRU_CO\ : std_logic;
signal \FSM_TEST_inst_slow.counter_statZ0Z_1\ : std_logic;
signal \FSM_TEST_inst_slow.counter_stat_cry_3_THRU_CO\ : std_logic;
signal \FSM_TEST_inst_slow.counter_statZ0Z_4\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_statZ0Z_4\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_statZ0Z_5\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_statZ0Z_1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idle_cry_0_THRU_CO\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.N_126_1_i_cascade_\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.current_state_d_i_2\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idleZ0Z_7\ : std_logic;
signal \FSM_TEST_inst_slow.flag_input_regZ0\ : std_logic;
signal \FSM_TEST_inst_slow.counter_idleZ0Z_6\ : std_logic;
signal \FSM_TEST_inst_slow.current_state_RNO_3Z0Z_0\ : std_logic;
signal \FSM_TEST_inst_slow.current_state_RNO_4Z0Z_0_cascade_\ : std_logic;
signal \FSM_TEST_inst_slow.current_state_RNO_5Z0Z_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_2\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_3\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_4\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_5\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idle_cry_3_THRU_CO\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.flag_input_regZ0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.G_24_0_a4_1_4\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idle_cry_1_THRU_CO\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idle_cry_2_THRU_CO\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_4\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_3\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_5\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idlelde_2_cascade_\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1_cascade_\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.N_126_1_i\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_2\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.G_24_0_a4_1_5\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_6\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_19\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_20\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_21\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_22\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_23\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_86\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_84\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_85\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_82\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_83\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_12\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_52\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_7\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_8\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_9\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_53\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_10\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_11\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_54\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_55\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_50\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_51\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_5\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_6\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_56\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_69\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_68\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_67\ : std_logic;
signal \FSM_TEST_inst_slow.N_108_li_cascade_\ : std_logic;
signal \FSM_TEST_inst_slow.current_state_RNIR2L81_0Z0Z_1\ : std_logic;
signal \FSM_TEST_inst_slow.current_state_cnv_0_1\ : std_logic;
signal \FSM_TEST_inst_slow.N_108_li\ : std_logic;
signal \FSM_TEST_inst_slow.counter_dinZ0Z_3\ : std_logic;
signal \FSM_TEST_inst_slow.counter_dinZ0Z_2\ : std_logic;
signal \FSM_TEST_inst_slow.N_106_0\ : std_logic;
signal \FSM_TEST_inst_slow.current_state_RNO_8Z0Z_0_cascade_\ : std_logic;
signal \FSM_TEST_inst_slow.current_state_RNO_1Z0Z_0\ : std_logic;
signal \FSM_TEST_inst_slow.N_134\ : std_logic;
signal \FSM_TEST_inst_slow.current_state_RNO_2Z0Z_0_cascade_\ : std_logic;
signal s12_c : std_logic;
signal \config_register_latched_dec_inst.DYNCNF_1Z0Z_8\ : std_logic;
signal \config_register_latched_dec_inst.DYNCNF_1Z0Z_9\ : std_logic;
signal s13_c : std_logic;
signal \config_register_latched_dec_inst.DYNCNF_1Z0Z_0\ : std_logic;
signal \config_register_latched_dec_inst.DYNCNF_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_din_3_i_0_2_cascade_\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.G_24_0_o4_2_cascade_\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.G_24_0_a4_0_1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_statZ0Z_6\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_statZ0Z_3\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.G_24_0_a4_0_5\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.N_18_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.G_24_0_a4_0_6_cascade_\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.N_9_1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_4\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_5\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_2\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_3\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_13\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_14\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_18\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_24\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_78\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_77\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_25\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_26\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.CLK_uC_3Z0Z_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.CLK_uC_4Z0Z_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.CLK_uC_5Z0Z_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.CLK_uC_6Z0Z_0\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_57\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_60\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_58\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_59\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_61\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_66\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_64\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_65\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_62\ : std_logic;
signal \FSM_TEST_inst_slow.current_stateZ0Z_1\ : std_logic;
signal \FSM_TEST_inst_slow.bit_sequence_statZ0Z_63\ : std_logic;
signal \FSM_TEST_inst_slow.N_374_g\ : std_logic;
signal \counter_RNIFD27_2_cascade_\ : std_logic;
signal \N_3_0_cascade_\ : std_logic;
signal \N_2_0\ : std_logic;
signal \counter_RNISR1F_2\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_15\ : std_logic;
signal \clk_out_RNI3LEM_cascade_\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.N_100_li_cascade_\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5DZ0Z1_cascade_\ : std_logic;
signal \N_378_i\ : std_logic;
signal flag_signal : std_logic;
signal mosi_fast : std_logic;
signal mosi_slow : std_logic;
signal mosi_output_c : std_logic;
signal \config_register_latched_dec_inst.DYNCNF_1Z0Z_10\ : std_logic;
signal s14_c : std_logic;
signal \config_register_latched_dec_inst.N_378_i_i\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.N_101_0\ : std_logic;
signal \config_register_latched_dec_inst.DYNSRZ0Z_10\ : std_logic;
signal miso_input_c : std_logic;
signal \config_register_latched_dec_inst.DYNSRZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_10\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_6\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_7\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_8\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_9\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_11\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_12\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.current_state_fast_RNI78E11Z0Z_1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_27\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_28\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_59\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_76\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_54\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.CLK_uC_2Z0Z_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.CLK_uC_6bZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.CLK_uCZ0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5DZ0Z1\ : std_logic;
signal \N_3_0\ : std_logic;
signal \N_4_0\ : std_logic;
signal \CLK_uC_6c_0\ : std_logic;
signal clk_output_c : std_logic;
signal \FSM_TEST_inst_slow.current_state_RNI9C3K2Z0Z_1\ : std_logic;
signal \FSM_TEST_inst_slow.current_state_d_i_2\ : std_logic;
signal \FSM_TEST_inst_slow.counter_stat_cry_4_THRU_CO\ : std_logic;
signal \FSM_TEST_inst_slow.counter_statZ0Z_5\ : std_logic;
signal \divisor_inst_2.counterZ0Z_1\ : std_logic;
signal \divisor_inst_2.counterZ0Z_0\ : std_logic;
signal \divisor_inst_2.counterZ0Z_2\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.aux_selection_fast_0\ : std_logic;
signal \FSM_TEST_inst_slow.current_stateZ1Z_0\ : std_logic;
signal \counter_RNIFD27_2\ : std_logic;
signal clk_continuous_slow : std_logic;
signal \FSM_TEST_inst_slow.aux_selection_slow_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.current_state_fast_fastZ0Z_1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.current_state_fast_1_repZ0Z1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.current_state_fastZ0Z_1\ : std_logic;
signal \FSM_TEST_inst_slow.CLK_uC_6kZ0Z_0\ : std_logic;
signal \CLK_uC_6l_0\ : std_logic;
signal \config_register_latched_dec_inst.DYNSRZ0Z_3\ : std_logic;
signal \config_register_latched_dec_inst.DYNSRZ0Z_4\ : std_logic;
signal \config_register_latched_dec_inst.DYNSRZ0Z_1\ : std_logic;
signal \config_register_latched_dec_inst.DYNSRZ0Z_2\ : std_logic;
signal \config_register_latched_dec_inst.DYNSRZ0Z_7\ : std_logic;
signal \config_register_latched_dec_inst.DYNSRZ0Z_5\ : std_logic;
signal \config_register_latched_dec_inst.DYNSRZ0Z_6\ : std_logic;
signal \config_register_latched_dec_inst.DYNSRZ0Z_8\ : std_logic;
signal \config_register_latched_dec_inst.DYNSRZ0Z_9\ : std_logic;
signal \flag_output_0_ret_RNI1E8NZ0Z2\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_51\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_52\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_53\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_31\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_50\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_29\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_30\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_75\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_60\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_58\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_7\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_8\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_9\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_57\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_79\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_55\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_56\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_83\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_87\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_84\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_85\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_86\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_82\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_65\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_35\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_80\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_81\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_32\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_39\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_46\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_47\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_40\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_48\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_49\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_33\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_34\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_10\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_74\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_13\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_14\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_15\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_16\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_17\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_11\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_12\ : std_logic;
signal \config_register_latched_dec_inst.STATSRZ0Z_0\ : std_logic;
signal \config_register_latched_dec_inst.STATCNF_1Z0Z_0\ : std_logic;
signal sel_output_c : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_2\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_dinZ1Z_1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_3\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_66\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_67\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_45\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_38\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_36\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_37\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_43\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_44\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_64\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_63\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_61\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_62\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_68\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_41\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_42\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_69\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_70\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_71\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_72\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_73\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.N_256_g\ : std_logic;
signal \RST_N_c\ : std_logic;
signal \RST_N_c_i\ : std_logic;
signal divisor_inst_counter_0 : std_logic;
signal clk_continuous_fast : std_logic;
signal divisor_inst_counter_1 : std_logic;
signal \FSM_TEST_inst_RAPIDA.N_100_li\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIKIU51Z0Z_1\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z2\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.N_123_0\ : std_logic;
signal \clk_out_RNI3LEM\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.current_stateZ0Z_0\ : std_logic;
signal \FSM_TEST_inst_RAPIDA.current_stateZ0Z_1\ : std_logic;
signal clk_pll_1 : std_logic;
signal \RST_N_c_i_g\ : std_logic;
signal \config_register_latched_dec_inst.STATCNF_0\ : std_logic;
signal \STATCNF_i_0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal xor_out_stat_wire : std_logic;
signal clk_output_wire : std_logic;
signal s13_wire : std_logic;
signal sel_output_wire : std_logic;
signal xor_out_dyn_wire : std_logic;
signal s12_wire : std_logic;
signal miso_input_wire : std_logic;
signal \RST_N_wire\ : std_logic;
signal mosi_output_wire : std_logic;
signal s14_wire : std_logic;
signal \top_pll_inst.top_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK_wire\ <= CLK;
    xor_out_stat <= xor_out_stat_wire;
    clk_output <= clk_output_wire;
    s13 <= s13_wire;
    sel_output <= sel_output_wire;
    xor_out_dyn <= xor_out_dyn_wire;
    s12 <= s12_wire;
    miso_input_wire <= miso_input;
    \RST_N_wire\ <= RST_N;
    mosi_output <= mosi_output_wire;
    s14 <= s14_wire;
    \top_pll_inst.top_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \top_pll_inst.top_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__4904\,
            RESETB => \N__12104\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \top_pll_inst.top_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_pll_1
        );

    \CLK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12279\,
            DIN => \N__12278\,
            DOUT => \N__12277\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12279\,
            PADOUT => \N__12278\,
            PADIN => \N__12277\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \xor_out_stat_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12270\,
            DIN => \N__12269\,
            DOUT => \N__12268\,
            PACKAGEPIN => xor_out_stat_wire
        );

    \xor_out_stat_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12270\,
            PADOUT => \N__12269\,
            PADIN => \N__12268\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10442\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12261\,
            DIN => \N__12260\,
            DOUT => \N__12259\,
            PACKAGEPIN => clk_output_wire
        );

    \clk_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12261\,
            PADOUT => \N__12260\,
            PADIN => \N__12259\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8303\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s13_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12252\,
            DIN => \N__12251\,
            DOUT => \N__12250\,
            PACKAGEPIN => s13_wire
        );

    \s13_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12252\,
            PADOUT => \N__12251\,
            PADIN => \N__12250\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6812\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sel_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12243\,
            DIN => \N__12242\,
            DOUT => \N__12241\,
            PACKAGEPIN => sel_output_wire
        );

    \sel_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12243\,
            PADOUT => \N__12242\,
            PADIN => \N__12241\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10112\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \xor_out_dyn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12234\,
            DIN => \N__12233\,
            DOUT => \N__12232\,
            PACKAGEPIN => xor_out_dyn_wire
        );

    \xor_out_dyn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12234\,
            PADOUT => \N__12233\,
            PADIN => \N__12232\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4958\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s12_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12225\,
            DIN => \N__12224\,
            DOUT => \N__12223\,
            PACKAGEPIN => s12_wire
        );

    \s12_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12225\,
            PADOUT => \N__12224\,
            PADIN => \N__12223\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6854\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \miso_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12216\,
            DIN => \N__12215\,
            DOUT => \N__12214\,
            PACKAGEPIN => miso_input_wire
        );

    \miso_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12216\,
            PADOUT => \N__12215\,
            PADIN => \N__12214\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => miso_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RST_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12207\,
            DIN => \N__12206\,
            DOUT => \N__12205\,
            PACKAGEPIN => \RST_N_wire\
        );

    \RST_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12207\,
            PADOUT => \N__12206\,
            PADIN => \N__12205\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RST_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \mosi_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12198\,
            DIN => \N__12197\,
            DOUT => \N__12196\,
            PACKAGEPIN => mosi_output_wire
        );

    \mosi_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12198\,
            PADOUT => \N__12197\,
            PADIN => \N__12196\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8027\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s14_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12189\,
            DIN => \N__12188\,
            DOUT => \N__12187\,
            PACKAGEPIN => s14_wire
        );

    \s14_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12189\,
            PADOUT => \N__12188\,
            PADIN => \N__12187\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7985\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2841\ : InMux
    port map (
            O => \N__12170\,
            I => \N__12167\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__12167\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_71\
        );

    \I__2839\ : InMux
    port map (
            O => \N__12164\,
            I => \N__12161\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__12161\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_72\
        );

    \I__2837\ : InMux
    port map (
            O => \N__12158\,
            I => \N__12155\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__12155\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_73\
        );

    \I__2835\ : CEMux
    port map (
            O => \N__12152\,
            I => \N__12110\
        );

    \I__2834\ : CEMux
    port map (
            O => \N__12151\,
            I => \N__12110\
        );

    \I__2833\ : CEMux
    port map (
            O => \N__12150\,
            I => \N__12110\
        );

    \I__2832\ : CEMux
    port map (
            O => \N__12149\,
            I => \N__12110\
        );

    \I__2831\ : CEMux
    port map (
            O => \N__12148\,
            I => \N__12110\
        );

    \I__2830\ : CEMux
    port map (
            O => \N__12147\,
            I => \N__12110\
        );

    \I__2829\ : CEMux
    port map (
            O => \N__12146\,
            I => \N__12110\
        );

    \I__2828\ : CEMux
    port map (
            O => \N__12145\,
            I => \N__12110\
        );

    \I__2827\ : CEMux
    port map (
            O => \N__12144\,
            I => \N__12110\
        );

    \I__2826\ : CEMux
    port map (
            O => \N__12143\,
            I => \N__12110\
        );

    \I__2825\ : CEMux
    port map (
            O => \N__12142\,
            I => \N__12110\
        );

    \I__2824\ : CEMux
    port map (
            O => \N__12141\,
            I => \N__12110\
        );

    \I__2823\ : CEMux
    port map (
            O => \N__12140\,
            I => \N__12110\
        );

    \I__2822\ : CEMux
    port map (
            O => \N__12139\,
            I => \N__12110\
        );

    \I__2821\ : GlobalMux
    port map (
            O => \N__12110\,
            I => \N__12107\
        );

    \I__2820\ : gio2CtrlBuf
    port map (
            O => \N__12107\,
            I => \FSM_TEST_inst_RAPIDA.N_256_g\
        );

    \I__2819\ : IoInMux
    port map (
            O => \N__12104\,
            I => \N__12101\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__12101\,
            I => \N__12098\
        );

    \I__2817\ : IoSpan4Mux
    port map (
            O => \N__12098\,
            I => \N__12092\
        );

    \I__2816\ : InMux
    port map (
            O => \N__12097\,
            I => \N__12089\
        );

    \I__2815\ : InMux
    port map (
            O => \N__12096\,
            I => \N__12084\
        );

    \I__2814\ : InMux
    port map (
            O => \N__12095\,
            I => \N__12084\
        );

    \I__2813\ : Span4Mux_s3_v
    port map (
            O => \N__12092\,
            I => \N__12078\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__12089\,
            I => \N__12075\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__12084\,
            I => \N__12072\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__12083\,
            I => \N__12067\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__12082\,
            I => \N__12064\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__12081\,
            I => \N__12059\
        );

    \I__2807\ : Sp12to4
    port map (
            O => \N__12078\,
            I => \N__12056\
        );

    \I__2806\ : Span4Mux_v
    port map (
            O => \N__12075\,
            I => \N__12053\
        );

    \I__2805\ : Span4Mux_v
    port map (
            O => \N__12072\,
            I => \N__12050\
        );

    \I__2804\ : InMux
    port map (
            O => \N__12071\,
            I => \N__12035\
        );

    \I__2803\ : InMux
    port map (
            O => \N__12070\,
            I => \N__12035\
        );

    \I__2802\ : InMux
    port map (
            O => \N__12067\,
            I => \N__12035\
        );

    \I__2801\ : InMux
    port map (
            O => \N__12064\,
            I => \N__12035\
        );

    \I__2800\ : InMux
    port map (
            O => \N__12063\,
            I => \N__12035\
        );

    \I__2799\ : InMux
    port map (
            O => \N__12062\,
            I => \N__12035\
        );

    \I__2798\ : InMux
    port map (
            O => \N__12059\,
            I => \N__12035\
        );

    \I__2797\ : Span12Mux_v
    port map (
            O => \N__12056\,
            I => \N__12025\
        );

    \I__2796\ : Sp12to4
    port map (
            O => \N__12053\,
            I => \N__12025\
        );

    \I__2795\ : Sp12to4
    port map (
            O => \N__12050\,
            I => \N__12025\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__12035\,
            I => \N__12025\
        );

    \I__2793\ : InMux
    port map (
            O => \N__12034\,
            I => \N__12022\
        );

    \I__2792\ : Span12Mux_h
    port map (
            O => \N__12025\,
            I => \N__12019\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__12022\,
            I => \N__12016\
        );

    \I__2790\ : Span12Mux_v
    port map (
            O => \N__12019\,
            I => \N__12011\
        );

    \I__2789\ : Span12Mux_h
    port map (
            O => \N__12016\,
            I => \N__12011\
        );

    \I__2788\ : Odrv12
    port map (
            O => \N__12011\,
            I => \RST_N_c\
        );

    \I__2787\ : IoInMux
    port map (
            O => \N__12008\,
            I => \N__12005\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__12005\,
            I => \N__12002\
        );

    \I__2785\ : Odrv12
    port map (
            O => \N__12002\,
            I => \RST_N_c_i\
        );

    \I__2784\ : InMux
    port map (
            O => \N__11999\,
            I => \N__11993\
        );

    \I__2783\ : InMux
    port map (
            O => \N__11998\,
            I => \N__11985\
        );

    \I__2782\ : InMux
    port map (
            O => \N__11997\,
            I => \N__11985\
        );

    \I__2781\ : InMux
    port map (
            O => \N__11996\,
            I => \N__11985\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__11993\,
            I => \N__11982\
        );

    \I__2779\ : InMux
    port map (
            O => \N__11992\,
            I => \N__11979\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__11985\,
            I => divisor_inst_counter_0
        );

    \I__2777\ : Odrv4
    port map (
            O => \N__11982\,
            I => divisor_inst_counter_0
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__11979\,
            I => divisor_inst_counter_0
        );

    \I__2775\ : InMux
    port map (
            O => \N__11972\,
            I => \N__11969\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__11969\,
            I => \N__11965\
        );

    \I__2773\ : InMux
    port map (
            O => \N__11968\,
            I => \N__11961\
        );

    \I__2772\ : Span4Mux_v
    port map (
            O => \N__11965\,
            I => \N__11957\
        );

    \I__2771\ : InMux
    port map (
            O => \N__11964\,
            I => \N__11954\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__11961\,
            I => \N__11951\
        );

    \I__2769\ : InMux
    port map (
            O => \N__11960\,
            I => \N__11948\
        );

    \I__2768\ : Odrv4
    port map (
            O => \N__11957\,
            I => clk_continuous_fast
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__11954\,
            I => clk_continuous_fast
        );

    \I__2766\ : Odrv4
    port map (
            O => \N__11951\,
            I => clk_continuous_fast
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__11948\,
            I => clk_continuous_fast
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__11939\,
            I => \N__11936\
        );

    \I__2763\ : InMux
    port map (
            O => \N__11936\,
            I => \N__11931\
        );

    \I__2762\ : InMux
    port map (
            O => \N__11935\,
            I => \N__11925\
        );

    \I__2761\ : InMux
    port map (
            O => \N__11934\,
            I => \N__11925\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__11931\,
            I => \N__11922\
        );

    \I__2759\ : InMux
    port map (
            O => \N__11930\,
            I => \N__11919\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__11925\,
            I => divisor_inst_counter_1
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__11922\,
            I => divisor_inst_counter_1
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__11919\,
            I => divisor_inst_counter_1
        );

    \I__2755\ : InMux
    port map (
            O => \N__11912\,
            I => \N__11905\
        );

    \I__2754\ : InMux
    port map (
            O => \N__11911\,
            I => \N__11902\
        );

    \I__2753\ : InMux
    port map (
            O => \N__11910\,
            I => \N__11895\
        );

    \I__2752\ : InMux
    port map (
            O => \N__11909\,
            I => \N__11895\
        );

    \I__2751\ : InMux
    port map (
            O => \N__11908\,
            I => \N__11895\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__11905\,
            I => \N__11892\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__11902\,
            I => \FSM_TEST_inst_RAPIDA.N_100_li\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__11895\,
            I => \FSM_TEST_inst_RAPIDA.N_100_li\
        );

    \I__2747\ : Odrv12
    port map (
            O => \N__11892\,
            I => \FSM_TEST_inst_RAPIDA.N_100_li\
        );

    \I__2746\ : IoInMux
    port map (
            O => \N__11885\,
            I => \N__11882\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__11882\,
            I => \N__11879\
        );

    \I__2744\ : Span12Mux_s5_v
    port map (
            O => \N__11879\,
            I => \N__11876\
        );

    \I__2743\ : Odrv12
    port map (
            O => \N__11876\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIKIU51Z0Z_1\
        );

    \I__2742\ : InMux
    port map (
            O => \N__11873\,
            I => \N__11854\
        );

    \I__2741\ : InMux
    port map (
            O => \N__11872\,
            I => \N__11854\
        );

    \I__2740\ : InMux
    port map (
            O => \N__11871\,
            I => \N__11854\
        );

    \I__2739\ : CascadeMux
    port map (
            O => \N__11870\,
            I => \N__11848\
        );

    \I__2738\ : InMux
    port map (
            O => \N__11869\,
            I => \N__11836\
        );

    \I__2737\ : InMux
    port map (
            O => \N__11868\,
            I => \N__11836\
        );

    \I__2736\ : InMux
    port map (
            O => \N__11867\,
            I => \N__11836\
        );

    \I__2735\ : InMux
    port map (
            O => \N__11866\,
            I => \N__11836\
        );

    \I__2734\ : InMux
    port map (
            O => \N__11865\,
            I => \N__11836\
        );

    \I__2733\ : InMux
    port map (
            O => \N__11864\,
            I => \N__11821\
        );

    \I__2732\ : InMux
    port map (
            O => \N__11863\,
            I => \N__11818\
        );

    \I__2731\ : InMux
    port map (
            O => \N__11862\,
            I => \N__11813\
        );

    \I__2730\ : InMux
    port map (
            O => \N__11861\,
            I => \N__11813\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__11854\,
            I => \N__11807\
        );

    \I__2728\ : InMux
    port map (
            O => \N__11853\,
            I => \N__11802\
        );

    \I__2727\ : InMux
    port map (
            O => \N__11852\,
            I => \N__11802\
        );

    \I__2726\ : InMux
    port map (
            O => \N__11851\,
            I => \N__11795\
        );

    \I__2725\ : InMux
    port map (
            O => \N__11848\,
            I => \N__11795\
        );

    \I__2724\ : InMux
    port map (
            O => \N__11847\,
            I => \N__11795\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__11836\,
            I => \N__11792\
        );

    \I__2722\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11781\
        );

    \I__2721\ : InMux
    port map (
            O => \N__11834\,
            I => \N__11781\
        );

    \I__2720\ : InMux
    port map (
            O => \N__11833\,
            I => \N__11781\
        );

    \I__2719\ : InMux
    port map (
            O => \N__11832\,
            I => \N__11781\
        );

    \I__2718\ : InMux
    port map (
            O => \N__11831\,
            I => \N__11781\
        );

    \I__2717\ : InMux
    port map (
            O => \N__11830\,
            I => \N__11772\
        );

    \I__2716\ : InMux
    port map (
            O => \N__11829\,
            I => \N__11772\
        );

    \I__2715\ : InMux
    port map (
            O => \N__11828\,
            I => \N__11772\
        );

    \I__2714\ : InMux
    port map (
            O => \N__11827\,
            I => \N__11772\
        );

    \I__2713\ : InMux
    port map (
            O => \N__11826\,
            I => \N__11765\
        );

    \I__2712\ : InMux
    port map (
            O => \N__11825\,
            I => \N__11765\
        );

    \I__2711\ : InMux
    port map (
            O => \N__11824\,
            I => \N__11765\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__11821\,
            I => \N__11760\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__11818\,
            I => \N__11760\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__11813\,
            I => \N__11757\
        );

    \I__2707\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11750\
        );

    \I__2706\ : InMux
    port map (
            O => \N__11811\,
            I => \N__11750\
        );

    \I__2705\ : InMux
    port map (
            O => \N__11810\,
            I => \N__11750\
        );

    \I__2704\ : Span4Mux_h
    port map (
            O => \N__11807\,
            I => \N__11744\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__11802\,
            I => \N__11744\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__11795\,
            I => \N__11741\
        );

    \I__2701\ : Span4Mux_v
    port map (
            O => \N__11792\,
            I => \N__11736\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__11781\,
            I => \N__11736\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__11772\,
            I => \N__11731\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__11765\,
            I => \N__11731\
        );

    \I__2697\ : Span4Mux_v
    port map (
            O => \N__11760\,
            I => \N__11724\
        );

    \I__2696\ : Span4Mux_h
    port map (
            O => \N__11757\,
            I => \N__11724\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__11750\,
            I => \N__11724\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__11749\,
            I => \N__11720\
        );

    \I__2693\ : Span4Mux_v
    port map (
            O => \N__11744\,
            I => \N__11717\
        );

    \I__2692\ : Span4Mux_h
    port map (
            O => \N__11741\,
            I => \N__11712\
        );

    \I__2691\ : Span4Mux_h
    port map (
            O => \N__11736\,
            I => \N__11712\
        );

    \I__2690\ : Span4Mux_v
    port map (
            O => \N__11731\,
            I => \N__11707\
        );

    \I__2689\ : Span4Mux_h
    port map (
            O => \N__11724\,
            I => \N__11707\
        );

    \I__2688\ : InMux
    port map (
            O => \N__11723\,
            I => \N__11704\
        );

    \I__2687\ : InMux
    port map (
            O => \N__11720\,
            I => \N__11701\
        );

    \I__2686\ : Odrv4
    port map (
            O => \N__11717\,
            I => \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z2\
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__11712\,
            I => \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z2\
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__11707\,
            I => \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z2\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__11704\,
            I => \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z2\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__11701\,
            I => \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z2\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__11690\,
            I => \N__11686\
        );

    \I__2680\ : InMux
    port map (
            O => \N__11689\,
            I => \N__11675\
        );

    \I__2679\ : InMux
    port map (
            O => \N__11686\,
            I => \N__11675\
        );

    \I__2678\ : InMux
    port map (
            O => \N__11685\,
            I => \N__11675\
        );

    \I__2677\ : InMux
    port map (
            O => \N__11684\,
            I => \N__11675\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__11675\,
            I => \N__11672\
        );

    \I__2675\ : Span4Mux_h
    port map (
            O => \N__11672\,
            I => \N__11667\
        );

    \I__2674\ : InMux
    port map (
            O => \N__11671\,
            I => \N__11662\
        );

    \I__2673\ : InMux
    port map (
            O => \N__11670\,
            I => \N__11662\
        );

    \I__2672\ : Odrv4
    port map (
            O => \N__11667\,
            I => \FSM_TEST_inst_RAPIDA.N_123_0\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__11662\,
            I => \FSM_TEST_inst_RAPIDA.N_123_0\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__11657\,
            I => \N__11652\
        );

    \I__2669\ : InMux
    port map (
            O => \N__11656\,
            I => \N__11646\
        );

    \I__2668\ : InMux
    port map (
            O => \N__11655\,
            I => \N__11643\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11652\,
            I => \N__11639\
        );

    \I__2666\ : InMux
    port map (
            O => \N__11651\,
            I => \N__11636\
        );

    \I__2665\ : InMux
    port map (
            O => \N__11650\,
            I => \N__11633\
        );

    \I__2664\ : InMux
    port map (
            O => \N__11649\,
            I => \N__11630\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__11646\,
            I => \N__11625\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__11643\,
            I => \N__11625\
        );

    \I__2661\ : CEMux
    port map (
            O => \N__11642\,
            I => \N__11610\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__11639\,
            I => \N__11603\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__11636\,
            I => \N__11603\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__11633\,
            I => \N__11603\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__11630\,
            I => \N__11600\
        );

    \I__2656\ : Span4Mux_h
    port map (
            O => \N__11625\,
            I => \N__11595\
        );

    \I__2655\ : InMux
    port map (
            O => \N__11624\,
            I => \N__11584\
        );

    \I__2654\ : InMux
    port map (
            O => \N__11623\,
            I => \N__11584\
        );

    \I__2653\ : InMux
    port map (
            O => \N__11622\,
            I => \N__11584\
        );

    \I__2652\ : InMux
    port map (
            O => \N__11621\,
            I => \N__11584\
        );

    \I__2651\ : InMux
    port map (
            O => \N__11620\,
            I => \N__11584\
        );

    \I__2650\ : InMux
    port map (
            O => \N__11619\,
            I => \N__11581\
        );

    \I__2649\ : InMux
    port map (
            O => \N__11618\,
            I => \N__11578\
        );

    \I__2648\ : InMux
    port map (
            O => \N__11617\,
            I => \N__11567\
        );

    \I__2647\ : InMux
    port map (
            O => \N__11616\,
            I => \N__11567\
        );

    \I__2646\ : InMux
    port map (
            O => \N__11615\,
            I => \N__11567\
        );

    \I__2645\ : InMux
    port map (
            O => \N__11614\,
            I => \N__11567\
        );

    \I__2644\ : InMux
    port map (
            O => \N__11613\,
            I => \N__11567\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__11610\,
            I => \N__11562\
        );

    \I__2642\ : Span4Mux_v
    port map (
            O => \N__11603\,
            I => \N__11562\
        );

    \I__2641\ : Span4Mux_h
    port map (
            O => \N__11600\,
            I => \N__11559\
        );

    \I__2640\ : InMux
    port map (
            O => \N__11599\,
            I => \N__11556\
        );

    \I__2639\ : InMux
    port map (
            O => \N__11598\,
            I => \N__11553\
        );

    \I__2638\ : Odrv4
    port map (
            O => \N__11595\,
            I => \clk_out_RNI3LEM\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__11584\,
            I => \clk_out_RNI3LEM\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__11581\,
            I => \clk_out_RNI3LEM\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__11578\,
            I => \clk_out_RNI3LEM\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__11567\,
            I => \clk_out_RNI3LEM\
        );

    \I__2633\ : Odrv4
    port map (
            O => \N__11562\,
            I => \clk_out_RNI3LEM\
        );

    \I__2632\ : Odrv4
    port map (
            O => \N__11559\,
            I => \clk_out_RNI3LEM\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__11556\,
            I => \clk_out_RNI3LEM\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__11553\,
            I => \clk_out_RNI3LEM\
        );

    \I__2629\ : InMux
    port map (
            O => \N__11534\,
            I => \N__11490\
        );

    \I__2628\ : InMux
    port map (
            O => \N__11533\,
            I => \N__11439\
        );

    \I__2627\ : InMux
    port map (
            O => \N__11532\,
            I => \N__11439\
        );

    \I__2626\ : InMux
    port map (
            O => \N__11531\,
            I => \N__11439\
        );

    \I__2625\ : InMux
    port map (
            O => \N__11530\,
            I => \N__11439\
        );

    \I__2624\ : InMux
    port map (
            O => \N__11529\,
            I => \N__11439\
        );

    \I__2623\ : InMux
    port map (
            O => \N__11528\,
            I => \N__11439\
        );

    \I__2622\ : InMux
    port map (
            O => \N__11527\,
            I => \N__11439\
        );

    \I__2621\ : InMux
    port map (
            O => \N__11526\,
            I => \N__11426\
        );

    \I__2620\ : InMux
    port map (
            O => \N__11525\,
            I => \N__11426\
        );

    \I__2619\ : InMux
    port map (
            O => \N__11524\,
            I => \N__11426\
        );

    \I__2618\ : InMux
    port map (
            O => \N__11523\,
            I => \N__11426\
        );

    \I__2617\ : InMux
    port map (
            O => \N__11522\,
            I => \N__11426\
        );

    \I__2616\ : InMux
    port map (
            O => \N__11521\,
            I => \N__11426\
        );

    \I__2615\ : InMux
    port map (
            O => \N__11520\,
            I => \N__11409\
        );

    \I__2614\ : InMux
    port map (
            O => \N__11519\,
            I => \N__11409\
        );

    \I__2613\ : InMux
    port map (
            O => \N__11518\,
            I => \N__11409\
        );

    \I__2612\ : InMux
    port map (
            O => \N__11517\,
            I => \N__11409\
        );

    \I__2611\ : InMux
    port map (
            O => \N__11516\,
            I => \N__11409\
        );

    \I__2610\ : InMux
    port map (
            O => \N__11515\,
            I => \N__11409\
        );

    \I__2609\ : InMux
    port map (
            O => \N__11514\,
            I => \N__11409\
        );

    \I__2608\ : InMux
    port map (
            O => \N__11513\,
            I => \N__11409\
        );

    \I__2607\ : InMux
    port map (
            O => \N__11512\,
            I => \N__11402\
        );

    \I__2606\ : InMux
    port map (
            O => \N__11511\,
            I => \N__11402\
        );

    \I__2605\ : InMux
    port map (
            O => \N__11510\,
            I => \N__11402\
        );

    \I__2604\ : InMux
    port map (
            O => \N__11509\,
            I => \N__11385\
        );

    \I__2603\ : InMux
    port map (
            O => \N__11508\,
            I => \N__11385\
        );

    \I__2602\ : InMux
    port map (
            O => \N__11507\,
            I => \N__11385\
        );

    \I__2601\ : InMux
    port map (
            O => \N__11506\,
            I => \N__11385\
        );

    \I__2600\ : InMux
    port map (
            O => \N__11505\,
            I => \N__11385\
        );

    \I__2599\ : InMux
    port map (
            O => \N__11504\,
            I => \N__11385\
        );

    \I__2598\ : InMux
    port map (
            O => \N__11503\,
            I => \N__11385\
        );

    \I__2597\ : InMux
    port map (
            O => \N__11502\,
            I => \N__11385\
        );

    \I__2596\ : InMux
    port map (
            O => \N__11501\,
            I => \N__11370\
        );

    \I__2595\ : InMux
    port map (
            O => \N__11500\,
            I => \N__11370\
        );

    \I__2594\ : InMux
    port map (
            O => \N__11499\,
            I => \N__11370\
        );

    \I__2593\ : InMux
    port map (
            O => \N__11498\,
            I => \N__11370\
        );

    \I__2592\ : InMux
    port map (
            O => \N__11497\,
            I => \N__11370\
        );

    \I__2591\ : InMux
    port map (
            O => \N__11496\,
            I => \N__11370\
        );

    \I__2590\ : InMux
    port map (
            O => \N__11495\,
            I => \N__11370\
        );

    \I__2589\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11361\
        );

    \I__2588\ : InMux
    port map (
            O => \N__11493\,
            I => \N__11361\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__11490\,
            I => \N__11358\
        );

    \I__2586\ : InMux
    port map (
            O => \N__11489\,
            I => \N__11343\
        );

    \I__2585\ : InMux
    port map (
            O => \N__11488\,
            I => \N__11343\
        );

    \I__2584\ : InMux
    port map (
            O => \N__11487\,
            I => \N__11343\
        );

    \I__2583\ : InMux
    port map (
            O => \N__11486\,
            I => \N__11343\
        );

    \I__2582\ : InMux
    port map (
            O => \N__11485\,
            I => \N__11343\
        );

    \I__2581\ : InMux
    port map (
            O => \N__11484\,
            I => \N__11343\
        );

    \I__2580\ : InMux
    port map (
            O => \N__11483\,
            I => \N__11343\
        );

    \I__2579\ : InMux
    port map (
            O => \N__11482\,
            I => \N__11330\
        );

    \I__2578\ : InMux
    port map (
            O => \N__11481\,
            I => \N__11330\
        );

    \I__2577\ : InMux
    port map (
            O => \N__11480\,
            I => \N__11330\
        );

    \I__2576\ : InMux
    port map (
            O => \N__11479\,
            I => \N__11330\
        );

    \I__2575\ : InMux
    port map (
            O => \N__11478\,
            I => \N__11330\
        );

    \I__2574\ : InMux
    port map (
            O => \N__11477\,
            I => \N__11330\
        );

    \I__2573\ : InMux
    port map (
            O => \N__11476\,
            I => \N__11323\
        );

    \I__2572\ : InMux
    port map (
            O => \N__11475\,
            I => \N__11323\
        );

    \I__2571\ : InMux
    port map (
            O => \N__11474\,
            I => \N__11323\
        );

    \I__2570\ : InMux
    port map (
            O => \N__11473\,
            I => \N__11308\
        );

    \I__2569\ : InMux
    port map (
            O => \N__11472\,
            I => \N__11308\
        );

    \I__2568\ : InMux
    port map (
            O => \N__11471\,
            I => \N__11308\
        );

    \I__2567\ : InMux
    port map (
            O => \N__11470\,
            I => \N__11308\
        );

    \I__2566\ : InMux
    port map (
            O => \N__11469\,
            I => \N__11308\
        );

    \I__2565\ : InMux
    port map (
            O => \N__11468\,
            I => \N__11308\
        );

    \I__2564\ : InMux
    port map (
            O => \N__11467\,
            I => \N__11308\
        );

    \I__2563\ : InMux
    port map (
            O => \N__11466\,
            I => \N__11305\
        );

    \I__2562\ : InMux
    port map (
            O => \N__11465\,
            I => \N__11296\
        );

    \I__2561\ : InMux
    port map (
            O => \N__11464\,
            I => \N__11296\
        );

    \I__2560\ : InMux
    port map (
            O => \N__11463\,
            I => \N__11296\
        );

    \I__2559\ : InMux
    port map (
            O => \N__11462\,
            I => \N__11296\
        );

    \I__2558\ : InMux
    port map (
            O => \N__11461\,
            I => \N__11291\
        );

    \I__2557\ : InMux
    port map (
            O => \N__11460\,
            I => \N__11291\
        );

    \I__2556\ : InMux
    port map (
            O => \N__11459\,
            I => \N__11288\
        );

    \I__2555\ : InMux
    port map (
            O => \N__11458\,
            I => \N__11243\
        );

    \I__2554\ : InMux
    port map (
            O => \N__11457\,
            I => \N__11243\
        );

    \I__2553\ : InMux
    port map (
            O => \N__11456\,
            I => \N__11243\
        );

    \I__2552\ : InMux
    port map (
            O => \N__11455\,
            I => \N__11243\
        );

    \I__2551\ : InMux
    port map (
            O => \N__11454\,
            I => \N__11243\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__11439\,
            I => \N__11230\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__11426\,
            I => \N__11230\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__11409\,
            I => \N__11230\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__11402\,
            I => \N__11230\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__11385\,
            I => \N__11230\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__11370\,
            I => \N__11230\
        );

    \I__2544\ : InMux
    port map (
            O => \N__11369\,
            I => \N__11221\
        );

    \I__2543\ : InMux
    port map (
            O => \N__11368\,
            I => \N__11221\
        );

    \I__2542\ : InMux
    port map (
            O => \N__11367\,
            I => \N__11221\
        );

    \I__2541\ : InMux
    port map (
            O => \N__11366\,
            I => \N__11221\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__11361\,
            I => \N__11214\
        );

    \I__2539\ : Span4Mux_v
    port map (
            O => \N__11358\,
            I => \N__11214\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__11343\,
            I => \N__11199\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__11330\,
            I => \N__11199\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__11323\,
            I => \N__11199\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__11308\,
            I => \N__11199\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__11305\,
            I => \N__11199\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__11296\,
            I => \N__11199\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__11291\,
            I => \N__11199\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__11288\,
            I => \N__11196\
        );

    \I__2530\ : InMux
    port map (
            O => \N__11287\,
            I => \N__11188\
        );

    \I__2529\ : InMux
    port map (
            O => \N__11286\,
            I => \N__11188\
        );

    \I__2528\ : InMux
    port map (
            O => \N__11285\,
            I => \N__11173\
        );

    \I__2527\ : InMux
    port map (
            O => \N__11284\,
            I => \N__11173\
        );

    \I__2526\ : InMux
    port map (
            O => \N__11283\,
            I => \N__11173\
        );

    \I__2525\ : InMux
    port map (
            O => \N__11282\,
            I => \N__11173\
        );

    \I__2524\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11173\
        );

    \I__2523\ : InMux
    port map (
            O => \N__11280\,
            I => \N__11173\
        );

    \I__2522\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11173\
        );

    \I__2521\ : InMux
    port map (
            O => \N__11278\,
            I => \N__11158\
        );

    \I__2520\ : InMux
    port map (
            O => \N__11277\,
            I => \N__11158\
        );

    \I__2519\ : InMux
    port map (
            O => \N__11276\,
            I => \N__11158\
        );

    \I__2518\ : InMux
    port map (
            O => \N__11275\,
            I => \N__11158\
        );

    \I__2517\ : InMux
    port map (
            O => \N__11274\,
            I => \N__11158\
        );

    \I__2516\ : InMux
    port map (
            O => \N__11273\,
            I => \N__11158\
        );

    \I__2515\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11158\
        );

    \I__2514\ : InMux
    port map (
            O => \N__11271\,
            I => \N__11153\
        );

    \I__2513\ : InMux
    port map (
            O => \N__11270\,
            I => \N__11153\
        );

    \I__2512\ : InMux
    port map (
            O => \N__11269\,
            I => \N__11150\
        );

    \I__2511\ : InMux
    port map (
            O => \N__11268\,
            I => \N__11140\
        );

    \I__2510\ : InMux
    port map (
            O => \N__11267\,
            I => \N__11140\
        );

    \I__2509\ : InMux
    port map (
            O => \N__11266\,
            I => \N__11140\
        );

    \I__2508\ : InMux
    port map (
            O => \N__11265\,
            I => \N__11125\
        );

    \I__2507\ : InMux
    port map (
            O => \N__11264\,
            I => \N__11125\
        );

    \I__2506\ : InMux
    port map (
            O => \N__11263\,
            I => \N__11125\
        );

    \I__2505\ : InMux
    port map (
            O => \N__11262\,
            I => \N__11125\
        );

    \I__2504\ : InMux
    port map (
            O => \N__11261\,
            I => \N__11125\
        );

    \I__2503\ : InMux
    port map (
            O => \N__11260\,
            I => \N__11125\
        );

    \I__2502\ : InMux
    port map (
            O => \N__11259\,
            I => \N__11125\
        );

    \I__2501\ : InMux
    port map (
            O => \N__11258\,
            I => \N__11114\
        );

    \I__2500\ : InMux
    port map (
            O => \N__11257\,
            I => \N__11114\
        );

    \I__2499\ : InMux
    port map (
            O => \N__11256\,
            I => \N__11114\
        );

    \I__2498\ : InMux
    port map (
            O => \N__11255\,
            I => \N__11114\
        );

    \I__2497\ : InMux
    port map (
            O => \N__11254\,
            I => \N__11114\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__11243\,
            I => \N__11107\
        );

    \I__2495\ : Span4Mux_v
    port map (
            O => \N__11230\,
            I => \N__11107\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__11221\,
            I => \N__11107\
        );

    \I__2493\ : InMux
    port map (
            O => \N__11220\,
            I => \N__11104\
        );

    \I__2492\ : InMux
    port map (
            O => \N__11219\,
            I => \N__11101\
        );

    \I__2491\ : Span4Mux_h
    port map (
            O => \N__11214\,
            I => \N__11094\
        );

    \I__2490\ : Span4Mux_v
    port map (
            O => \N__11199\,
            I => \N__11094\
        );

    \I__2489\ : Span4Mux_v
    port map (
            O => \N__11196\,
            I => \N__11094\
        );

    \I__2488\ : InMux
    port map (
            O => \N__11195\,
            I => \N__11087\
        );

    \I__2487\ : InMux
    port map (
            O => \N__11194\,
            I => \N__11087\
        );

    \I__2486\ : InMux
    port map (
            O => \N__11193\,
            I => \N__11087\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__11188\,
            I => \N__11078\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__11173\,
            I => \N__11078\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__11158\,
            I => \N__11078\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__11153\,
            I => \N__11078\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__11150\,
            I => \N__11075\
        );

    \I__2480\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11068\
        );

    \I__2479\ : InMux
    port map (
            O => \N__11148\,
            I => \N__11068\
        );

    \I__2478\ : InMux
    port map (
            O => \N__11147\,
            I => \N__11068\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__11140\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_0\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__11125\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_0\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__11114\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_0\
        );

    \I__2474\ : Odrv4
    port map (
            O => \N__11107\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_0\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__11104\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_0\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__11101\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_0\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__11094\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_0\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__11087\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_0\
        );

    \I__2469\ : Odrv4
    port map (
            O => \N__11078\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_0\
        );

    \I__2468\ : Odrv4
    port map (
            O => \N__11075\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_0\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__11068\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_0\
        );

    \I__2466\ : InMux
    port map (
            O => \N__11045\,
            I => \N__11034\
        );

    \I__2465\ : InMux
    port map (
            O => \N__11044\,
            I => \N__11034\
        );

    \I__2464\ : InMux
    port map (
            O => \N__11043\,
            I => \N__11011\
        );

    \I__2463\ : InMux
    port map (
            O => \N__11042\,
            I => \N__11011\
        );

    \I__2462\ : InMux
    port map (
            O => \N__11041\,
            I => \N__11011\
        );

    \I__2461\ : InMux
    port map (
            O => \N__11040\,
            I => \N__11011\
        );

    \I__2460\ : InMux
    port map (
            O => \N__11039\,
            I => \N__11011\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__11034\,
            I => \N__11008\
        );

    \I__2458\ : InMux
    port map (
            O => \N__11033\,
            I => \N__11005\
        );

    \I__2457\ : InMux
    port map (
            O => \N__11032\,
            I => \N__10996\
        );

    \I__2456\ : InMux
    port map (
            O => \N__11031\,
            I => \N__10989\
        );

    \I__2455\ : InMux
    port map (
            O => \N__11030\,
            I => \N__10989\
        );

    \I__2454\ : InMux
    port map (
            O => \N__11029\,
            I => \N__10989\
        );

    \I__2453\ : InMux
    port map (
            O => \N__11028\,
            I => \N__10982\
        );

    \I__2452\ : InMux
    port map (
            O => \N__11027\,
            I => \N__10982\
        );

    \I__2451\ : InMux
    port map (
            O => \N__11026\,
            I => \N__10982\
        );

    \I__2450\ : InMux
    port map (
            O => \N__11025\,
            I => \N__10973\
        );

    \I__2449\ : InMux
    port map (
            O => \N__11024\,
            I => \N__10973\
        );

    \I__2448\ : InMux
    port map (
            O => \N__11023\,
            I => \N__10973\
        );

    \I__2447\ : InMux
    port map (
            O => \N__11022\,
            I => \N__10973\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__11011\,
            I => \N__10964\
        );

    \I__2445\ : Span4Mux_h
    port map (
            O => \N__11008\,
            I => \N__10959\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__11005\,
            I => \N__10959\
        );

    \I__2443\ : InMux
    port map (
            O => \N__11004\,
            I => \N__10952\
        );

    \I__2442\ : InMux
    port map (
            O => \N__11003\,
            I => \N__10952\
        );

    \I__2441\ : InMux
    port map (
            O => \N__11002\,
            I => \N__10952\
        );

    \I__2440\ : InMux
    port map (
            O => \N__11001\,
            I => \N__10945\
        );

    \I__2439\ : InMux
    port map (
            O => \N__11000\,
            I => \N__10945\
        );

    \I__2438\ : InMux
    port map (
            O => \N__10999\,
            I => \N__10945\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__10996\,
            I => \N__10934\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__10989\,
            I => \N__10934\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__10982\,
            I => \N__10934\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__10973\,
            I => \N__10934\
        );

    \I__2433\ : InMux
    port map (
            O => \N__10972\,
            I => \N__10923\
        );

    \I__2432\ : InMux
    port map (
            O => \N__10971\,
            I => \N__10923\
        );

    \I__2431\ : InMux
    port map (
            O => \N__10970\,
            I => \N__10923\
        );

    \I__2430\ : InMux
    port map (
            O => \N__10969\,
            I => \N__10923\
        );

    \I__2429\ : InMux
    port map (
            O => \N__10968\,
            I => \N__10923\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__10967\,
            I => \N__10920\
        );

    \I__2427\ : Span4Mux_h
    port map (
            O => \N__10964\,
            I => \N__10911\
        );

    \I__2426\ : Span4Mux_h
    port map (
            O => \N__10959\,
            I => \N__10911\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__10952\,
            I => \N__10911\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__10945\,
            I => \N__10911\
        );

    \I__2423\ : InMux
    port map (
            O => \N__10944\,
            I => \N__10906\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10943\,
            I => \N__10906\
        );

    \I__2421\ : Span4Mux_v
    port map (
            O => \N__10934\,
            I => \N__10901\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__10923\,
            I => \N__10901\
        );

    \I__2419\ : InMux
    port map (
            O => \N__10920\,
            I => \N__10898\
        );

    \I__2418\ : Odrv4
    port map (
            O => \N__10911\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_1\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__10906\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_1\
        );

    \I__2416\ : Odrv4
    port map (
            O => \N__10901\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_1\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__10898\,
            I => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_1\
        );

    \I__2414\ : ClkMux
    port map (
            O => \N__10889\,
            I => \N__10676\
        );

    \I__2413\ : ClkMux
    port map (
            O => \N__10888\,
            I => \N__10676\
        );

    \I__2412\ : ClkMux
    port map (
            O => \N__10887\,
            I => \N__10676\
        );

    \I__2411\ : ClkMux
    port map (
            O => \N__10886\,
            I => \N__10676\
        );

    \I__2410\ : ClkMux
    port map (
            O => \N__10885\,
            I => \N__10676\
        );

    \I__2409\ : ClkMux
    port map (
            O => \N__10884\,
            I => \N__10676\
        );

    \I__2408\ : ClkMux
    port map (
            O => \N__10883\,
            I => \N__10676\
        );

    \I__2407\ : ClkMux
    port map (
            O => \N__10882\,
            I => \N__10676\
        );

    \I__2406\ : ClkMux
    port map (
            O => \N__10881\,
            I => \N__10676\
        );

    \I__2405\ : ClkMux
    port map (
            O => \N__10880\,
            I => \N__10676\
        );

    \I__2404\ : ClkMux
    port map (
            O => \N__10879\,
            I => \N__10676\
        );

    \I__2403\ : ClkMux
    port map (
            O => \N__10878\,
            I => \N__10676\
        );

    \I__2402\ : ClkMux
    port map (
            O => \N__10877\,
            I => \N__10676\
        );

    \I__2401\ : ClkMux
    port map (
            O => \N__10876\,
            I => \N__10676\
        );

    \I__2400\ : ClkMux
    port map (
            O => \N__10875\,
            I => \N__10676\
        );

    \I__2399\ : ClkMux
    port map (
            O => \N__10874\,
            I => \N__10676\
        );

    \I__2398\ : ClkMux
    port map (
            O => \N__10873\,
            I => \N__10676\
        );

    \I__2397\ : ClkMux
    port map (
            O => \N__10872\,
            I => \N__10676\
        );

    \I__2396\ : ClkMux
    port map (
            O => \N__10871\,
            I => \N__10676\
        );

    \I__2395\ : ClkMux
    port map (
            O => \N__10870\,
            I => \N__10676\
        );

    \I__2394\ : ClkMux
    port map (
            O => \N__10869\,
            I => \N__10676\
        );

    \I__2393\ : ClkMux
    port map (
            O => \N__10868\,
            I => \N__10676\
        );

    \I__2392\ : ClkMux
    port map (
            O => \N__10867\,
            I => \N__10676\
        );

    \I__2391\ : ClkMux
    port map (
            O => \N__10866\,
            I => \N__10676\
        );

    \I__2390\ : ClkMux
    port map (
            O => \N__10865\,
            I => \N__10676\
        );

    \I__2389\ : ClkMux
    port map (
            O => \N__10864\,
            I => \N__10676\
        );

    \I__2388\ : ClkMux
    port map (
            O => \N__10863\,
            I => \N__10676\
        );

    \I__2387\ : ClkMux
    port map (
            O => \N__10862\,
            I => \N__10676\
        );

    \I__2386\ : ClkMux
    port map (
            O => \N__10861\,
            I => \N__10676\
        );

    \I__2385\ : ClkMux
    port map (
            O => \N__10860\,
            I => \N__10676\
        );

    \I__2384\ : ClkMux
    port map (
            O => \N__10859\,
            I => \N__10676\
        );

    \I__2383\ : ClkMux
    port map (
            O => \N__10858\,
            I => \N__10676\
        );

    \I__2382\ : ClkMux
    port map (
            O => \N__10857\,
            I => \N__10676\
        );

    \I__2381\ : ClkMux
    port map (
            O => \N__10856\,
            I => \N__10676\
        );

    \I__2380\ : ClkMux
    port map (
            O => \N__10855\,
            I => \N__10676\
        );

    \I__2379\ : ClkMux
    port map (
            O => \N__10854\,
            I => \N__10676\
        );

    \I__2378\ : ClkMux
    port map (
            O => \N__10853\,
            I => \N__10676\
        );

    \I__2377\ : ClkMux
    port map (
            O => \N__10852\,
            I => \N__10676\
        );

    \I__2376\ : ClkMux
    port map (
            O => \N__10851\,
            I => \N__10676\
        );

    \I__2375\ : ClkMux
    port map (
            O => \N__10850\,
            I => \N__10676\
        );

    \I__2374\ : ClkMux
    port map (
            O => \N__10849\,
            I => \N__10676\
        );

    \I__2373\ : ClkMux
    port map (
            O => \N__10848\,
            I => \N__10676\
        );

    \I__2372\ : ClkMux
    port map (
            O => \N__10847\,
            I => \N__10676\
        );

    \I__2371\ : ClkMux
    port map (
            O => \N__10846\,
            I => \N__10676\
        );

    \I__2370\ : ClkMux
    port map (
            O => \N__10845\,
            I => \N__10676\
        );

    \I__2369\ : ClkMux
    port map (
            O => \N__10844\,
            I => \N__10676\
        );

    \I__2368\ : ClkMux
    port map (
            O => \N__10843\,
            I => \N__10676\
        );

    \I__2367\ : ClkMux
    port map (
            O => \N__10842\,
            I => \N__10676\
        );

    \I__2366\ : ClkMux
    port map (
            O => \N__10841\,
            I => \N__10676\
        );

    \I__2365\ : ClkMux
    port map (
            O => \N__10840\,
            I => \N__10676\
        );

    \I__2364\ : ClkMux
    port map (
            O => \N__10839\,
            I => \N__10676\
        );

    \I__2363\ : ClkMux
    port map (
            O => \N__10838\,
            I => \N__10676\
        );

    \I__2362\ : ClkMux
    port map (
            O => \N__10837\,
            I => \N__10676\
        );

    \I__2361\ : ClkMux
    port map (
            O => \N__10836\,
            I => \N__10676\
        );

    \I__2360\ : ClkMux
    port map (
            O => \N__10835\,
            I => \N__10676\
        );

    \I__2359\ : ClkMux
    port map (
            O => \N__10834\,
            I => \N__10676\
        );

    \I__2358\ : ClkMux
    port map (
            O => \N__10833\,
            I => \N__10676\
        );

    \I__2357\ : ClkMux
    port map (
            O => \N__10832\,
            I => \N__10676\
        );

    \I__2356\ : ClkMux
    port map (
            O => \N__10831\,
            I => \N__10676\
        );

    \I__2355\ : ClkMux
    port map (
            O => \N__10830\,
            I => \N__10676\
        );

    \I__2354\ : ClkMux
    port map (
            O => \N__10829\,
            I => \N__10676\
        );

    \I__2353\ : ClkMux
    port map (
            O => \N__10828\,
            I => \N__10676\
        );

    \I__2352\ : ClkMux
    port map (
            O => \N__10827\,
            I => \N__10676\
        );

    \I__2351\ : ClkMux
    port map (
            O => \N__10826\,
            I => \N__10676\
        );

    \I__2350\ : ClkMux
    port map (
            O => \N__10825\,
            I => \N__10676\
        );

    \I__2349\ : ClkMux
    port map (
            O => \N__10824\,
            I => \N__10676\
        );

    \I__2348\ : ClkMux
    port map (
            O => \N__10823\,
            I => \N__10676\
        );

    \I__2347\ : ClkMux
    port map (
            O => \N__10822\,
            I => \N__10676\
        );

    \I__2346\ : ClkMux
    port map (
            O => \N__10821\,
            I => \N__10676\
        );

    \I__2345\ : ClkMux
    port map (
            O => \N__10820\,
            I => \N__10676\
        );

    \I__2344\ : ClkMux
    port map (
            O => \N__10819\,
            I => \N__10676\
        );

    \I__2343\ : GlobalMux
    port map (
            O => \N__10676\,
            I => clk_pll_1
        );

    \I__2342\ : SRMux
    port map (
            O => \N__10673\,
            I => \N__10460\
        );

    \I__2341\ : SRMux
    port map (
            O => \N__10672\,
            I => \N__10460\
        );

    \I__2340\ : SRMux
    port map (
            O => \N__10671\,
            I => \N__10460\
        );

    \I__2339\ : SRMux
    port map (
            O => \N__10670\,
            I => \N__10460\
        );

    \I__2338\ : SRMux
    port map (
            O => \N__10669\,
            I => \N__10460\
        );

    \I__2337\ : SRMux
    port map (
            O => \N__10668\,
            I => \N__10460\
        );

    \I__2336\ : SRMux
    port map (
            O => \N__10667\,
            I => \N__10460\
        );

    \I__2335\ : SRMux
    port map (
            O => \N__10666\,
            I => \N__10460\
        );

    \I__2334\ : SRMux
    port map (
            O => \N__10665\,
            I => \N__10460\
        );

    \I__2333\ : SRMux
    port map (
            O => \N__10664\,
            I => \N__10460\
        );

    \I__2332\ : SRMux
    port map (
            O => \N__10663\,
            I => \N__10460\
        );

    \I__2331\ : SRMux
    port map (
            O => \N__10662\,
            I => \N__10460\
        );

    \I__2330\ : SRMux
    port map (
            O => \N__10661\,
            I => \N__10460\
        );

    \I__2329\ : SRMux
    port map (
            O => \N__10660\,
            I => \N__10460\
        );

    \I__2328\ : SRMux
    port map (
            O => \N__10659\,
            I => \N__10460\
        );

    \I__2327\ : SRMux
    port map (
            O => \N__10658\,
            I => \N__10460\
        );

    \I__2326\ : SRMux
    port map (
            O => \N__10657\,
            I => \N__10460\
        );

    \I__2325\ : SRMux
    port map (
            O => \N__10656\,
            I => \N__10460\
        );

    \I__2324\ : SRMux
    port map (
            O => \N__10655\,
            I => \N__10460\
        );

    \I__2323\ : SRMux
    port map (
            O => \N__10654\,
            I => \N__10460\
        );

    \I__2322\ : SRMux
    port map (
            O => \N__10653\,
            I => \N__10460\
        );

    \I__2321\ : SRMux
    port map (
            O => \N__10652\,
            I => \N__10460\
        );

    \I__2320\ : SRMux
    port map (
            O => \N__10651\,
            I => \N__10460\
        );

    \I__2319\ : SRMux
    port map (
            O => \N__10650\,
            I => \N__10460\
        );

    \I__2318\ : SRMux
    port map (
            O => \N__10649\,
            I => \N__10460\
        );

    \I__2317\ : SRMux
    port map (
            O => \N__10648\,
            I => \N__10460\
        );

    \I__2316\ : SRMux
    port map (
            O => \N__10647\,
            I => \N__10460\
        );

    \I__2315\ : SRMux
    port map (
            O => \N__10646\,
            I => \N__10460\
        );

    \I__2314\ : SRMux
    port map (
            O => \N__10645\,
            I => \N__10460\
        );

    \I__2313\ : SRMux
    port map (
            O => \N__10644\,
            I => \N__10460\
        );

    \I__2312\ : SRMux
    port map (
            O => \N__10643\,
            I => \N__10460\
        );

    \I__2311\ : SRMux
    port map (
            O => \N__10642\,
            I => \N__10460\
        );

    \I__2310\ : SRMux
    port map (
            O => \N__10641\,
            I => \N__10460\
        );

    \I__2309\ : SRMux
    port map (
            O => \N__10640\,
            I => \N__10460\
        );

    \I__2308\ : SRMux
    port map (
            O => \N__10639\,
            I => \N__10460\
        );

    \I__2307\ : SRMux
    port map (
            O => \N__10638\,
            I => \N__10460\
        );

    \I__2306\ : SRMux
    port map (
            O => \N__10637\,
            I => \N__10460\
        );

    \I__2305\ : SRMux
    port map (
            O => \N__10636\,
            I => \N__10460\
        );

    \I__2304\ : SRMux
    port map (
            O => \N__10635\,
            I => \N__10460\
        );

    \I__2303\ : SRMux
    port map (
            O => \N__10634\,
            I => \N__10460\
        );

    \I__2302\ : SRMux
    port map (
            O => \N__10633\,
            I => \N__10460\
        );

    \I__2301\ : SRMux
    port map (
            O => \N__10632\,
            I => \N__10460\
        );

    \I__2300\ : SRMux
    port map (
            O => \N__10631\,
            I => \N__10460\
        );

    \I__2299\ : SRMux
    port map (
            O => \N__10630\,
            I => \N__10460\
        );

    \I__2298\ : SRMux
    port map (
            O => \N__10629\,
            I => \N__10460\
        );

    \I__2297\ : SRMux
    port map (
            O => \N__10628\,
            I => \N__10460\
        );

    \I__2296\ : SRMux
    port map (
            O => \N__10627\,
            I => \N__10460\
        );

    \I__2295\ : SRMux
    port map (
            O => \N__10626\,
            I => \N__10460\
        );

    \I__2294\ : SRMux
    port map (
            O => \N__10625\,
            I => \N__10460\
        );

    \I__2293\ : SRMux
    port map (
            O => \N__10624\,
            I => \N__10460\
        );

    \I__2292\ : SRMux
    port map (
            O => \N__10623\,
            I => \N__10460\
        );

    \I__2291\ : SRMux
    port map (
            O => \N__10622\,
            I => \N__10460\
        );

    \I__2290\ : SRMux
    port map (
            O => \N__10621\,
            I => \N__10460\
        );

    \I__2289\ : SRMux
    port map (
            O => \N__10620\,
            I => \N__10460\
        );

    \I__2288\ : SRMux
    port map (
            O => \N__10619\,
            I => \N__10460\
        );

    \I__2287\ : SRMux
    port map (
            O => \N__10618\,
            I => \N__10460\
        );

    \I__2286\ : SRMux
    port map (
            O => \N__10617\,
            I => \N__10460\
        );

    \I__2285\ : SRMux
    port map (
            O => \N__10616\,
            I => \N__10460\
        );

    \I__2284\ : SRMux
    port map (
            O => \N__10615\,
            I => \N__10460\
        );

    \I__2283\ : SRMux
    port map (
            O => \N__10614\,
            I => \N__10460\
        );

    \I__2282\ : SRMux
    port map (
            O => \N__10613\,
            I => \N__10460\
        );

    \I__2281\ : SRMux
    port map (
            O => \N__10612\,
            I => \N__10460\
        );

    \I__2280\ : SRMux
    port map (
            O => \N__10611\,
            I => \N__10460\
        );

    \I__2279\ : SRMux
    port map (
            O => \N__10610\,
            I => \N__10460\
        );

    \I__2278\ : SRMux
    port map (
            O => \N__10609\,
            I => \N__10460\
        );

    \I__2277\ : SRMux
    port map (
            O => \N__10608\,
            I => \N__10460\
        );

    \I__2276\ : SRMux
    port map (
            O => \N__10607\,
            I => \N__10460\
        );

    \I__2275\ : SRMux
    port map (
            O => \N__10606\,
            I => \N__10460\
        );

    \I__2274\ : SRMux
    port map (
            O => \N__10605\,
            I => \N__10460\
        );

    \I__2273\ : SRMux
    port map (
            O => \N__10604\,
            I => \N__10460\
        );

    \I__2272\ : SRMux
    port map (
            O => \N__10603\,
            I => \N__10460\
        );

    \I__2271\ : GlobalMux
    port map (
            O => \N__10460\,
            I => \N__10457\
        );

    \I__2270\ : gio2CtrlBuf
    port map (
            O => \N__10457\,
            I => \RST_N_c_i_g\
        );

    \I__2269\ : InMux
    port map (
            O => \N__10454\,
            I => \N__10451\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__10451\,
            I => \N__10448\
        );

    \I__2267\ : Span4Mux_h
    port map (
            O => \N__10448\,
            I => \N__10445\
        );

    \I__2266\ : Odrv4
    port map (
            O => \N__10445\,
            I => \config_register_latched_dec_inst.STATCNF_0\
        );

    \I__2265\ : IoInMux
    port map (
            O => \N__10442\,
            I => \N__10439\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__10439\,
            I => \N__10436\
        );

    \I__2263\ : Span4Mux_s3_h
    port map (
            O => \N__10436\,
            I => \N__10433\
        );

    \I__2262\ : Span4Mux_h
    port map (
            O => \N__10433\,
            I => \N__10430\
        );

    \I__2261\ : Span4Mux_h
    port map (
            O => \N__10430\,
            I => \N__10427\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__10427\,
            I => \STATCNF_i_0\
        );

    \I__2259\ : InMux
    port map (
            O => \N__10424\,
            I => \N__10421\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__10421\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_37\
        );

    \I__2257\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10415\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__10415\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_43\
        );

    \I__2255\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10409\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__10409\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_44\
        );

    \I__2253\ : InMux
    port map (
            O => \N__10406\,
            I => \N__10403\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__10403\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_64\
        );

    \I__2251\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10397\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__10397\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_63\
        );

    \I__2249\ : InMux
    port map (
            O => \N__10394\,
            I => \N__10391\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__10391\,
            I => \N__10388\
        );

    \I__2247\ : Odrv4
    port map (
            O => \N__10388\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_61\
        );

    \I__2246\ : InMux
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__10382\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_62\
        );

    \I__2244\ : InMux
    port map (
            O => \N__10379\,
            I => \N__10376\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__10376\,
            I => \N__10373\
        );

    \I__2242\ : Odrv4
    port map (
            O => \N__10373\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_68\
        );

    \I__2241\ : InMux
    port map (
            O => \N__10370\,
            I => \N__10367\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__10367\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_41\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__10364\,
            I => \N__10361\
        );

    \I__2238\ : InMux
    port map (
            O => \N__10361\,
            I => \N__10358\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__10358\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_42\
        );

    \I__2236\ : InMux
    port map (
            O => \N__10355\,
            I => \N__10352\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__10352\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_69\
        );

    \I__2234\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10346\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__10346\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_70\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__10343\,
            I => \N__10321\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__10342\,
            I => \N__10318\
        );

    \I__2230\ : CascadeMux
    port map (
            O => \N__10341\,
            I => \N__10315\
        );

    \I__2229\ : InMux
    port map (
            O => \N__10340\,
            I => \N__10291\
        );

    \I__2228\ : InMux
    port map (
            O => \N__10339\,
            I => \N__10291\
        );

    \I__2227\ : InMux
    port map (
            O => \N__10338\,
            I => \N__10291\
        );

    \I__2226\ : InMux
    port map (
            O => \N__10337\,
            I => \N__10291\
        );

    \I__2225\ : InMux
    port map (
            O => \N__10336\,
            I => \N__10291\
        );

    \I__2224\ : InMux
    port map (
            O => \N__10335\,
            I => \N__10291\
        );

    \I__2223\ : InMux
    port map (
            O => \N__10334\,
            I => \N__10291\
        );

    \I__2222\ : InMux
    port map (
            O => \N__10333\,
            I => \N__10282\
        );

    \I__2221\ : InMux
    port map (
            O => \N__10332\,
            I => \N__10282\
        );

    \I__2220\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10282\
        );

    \I__2219\ : InMux
    port map (
            O => \N__10330\,
            I => \N__10282\
        );

    \I__2218\ : InMux
    port map (
            O => \N__10329\,
            I => \N__10279\
        );

    \I__2217\ : InMux
    port map (
            O => \N__10328\,
            I => \N__10272\
        );

    \I__2216\ : InMux
    port map (
            O => \N__10327\,
            I => \N__10272\
        );

    \I__2215\ : InMux
    port map (
            O => \N__10326\,
            I => \N__10272\
        );

    \I__2214\ : InMux
    port map (
            O => \N__10325\,
            I => \N__10267\
        );

    \I__2213\ : InMux
    port map (
            O => \N__10324\,
            I => \N__10267\
        );

    \I__2212\ : InMux
    port map (
            O => \N__10321\,
            I => \N__10260\
        );

    \I__2211\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10260\
        );

    \I__2210\ : InMux
    port map (
            O => \N__10315\,
            I => \N__10260\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__10314\,
            I => \N__10255\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__10313\,
            I => \N__10252\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__10312\,
            I => \N__10249\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__10311\,
            I => \N__10246\
        );

    \I__2205\ : InMux
    port map (
            O => \N__10310\,
            I => \N__10232\
        );

    \I__2204\ : InMux
    port map (
            O => \N__10309\,
            I => \N__10232\
        );

    \I__2203\ : InMux
    port map (
            O => \N__10308\,
            I => \N__10232\
        );

    \I__2202\ : InMux
    port map (
            O => \N__10307\,
            I => \N__10232\
        );

    \I__2201\ : InMux
    port map (
            O => \N__10306\,
            I => \N__10232\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__10291\,
            I => \N__10227\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__10282\,
            I => \N__10227\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__10279\,
            I => \N__10218\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__10272\,
            I => \N__10218\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__10267\,
            I => \N__10218\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__10260\,
            I => \N__10218\
        );

    \I__2194\ : InMux
    port map (
            O => \N__10259\,
            I => \N__10215\
        );

    \I__2193\ : InMux
    port map (
            O => \N__10258\,
            I => \N__10202\
        );

    \I__2192\ : InMux
    port map (
            O => \N__10255\,
            I => \N__10202\
        );

    \I__2191\ : InMux
    port map (
            O => \N__10252\,
            I => \N__10202\
        );

    \I__2190\ : InMux
    port map (
            O => \N__10249\,
            I => \N__10202\
        );

    \I__2189\ : InMux
    port map (
            O => \N__10246\,
            I => \N__10202\
        );

    \I__2188\ : InMux
    port map (
            O => \N__10245\,
            I => \N__10202\
        );

    \I__2187\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10199\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__10243\,
            I => \N__10196\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__10232\,
            I => \N__10193\
        );

    \I__2184\ : Span4Mux_v
    port map (
            O => \N__10227\,
            I => \N__10188\
        );

    \I__2183\ : Span4Mux_v
    port map (
            O => \N__10218\,
            I => \N__10188\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__10215\,
            I => \N__10181\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__10202\,
            I => \N__10181\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__10199\,
            I => \N__10181\
        );

    \I__2179\ : InMux
    port map (
            O => \N__10196\,
            I => \N__10178\
        );

    \I__2178\ : Odrv4
    port map (
            O => \N__10193\,
            I => \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z1\
        );

    \I__2177\ : Odrv4
    port map (
            O => \N__10188\,
            I => \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z1\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__10181\,
            I => \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z1\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__10178\,
            I => \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z1\
        );

    \I__2174\ : InMux
    port map (
            O => \N__10169\,
            I => \N__10166\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__10166\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_11\
        );

    \I__2172\ : InMux
    port map (
            O => \N__10163\,
            I => \N__10160\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__10160\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_12\
        );

    \I__2170\ : InMux
    port map (
            O => \N__10157\,
            I => \N__10154\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__10154\,
            I => \N__10150\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__10153\,
            I => \N__10146\
        );

    \I__2167\ : Span4Mux_v
    port map (
            O => \N__10150\,
            I => \N__10143\
        );

    \I__2166\ : InMux
    port map (
            O => \N__10149\,
            I => \N__10140\
        );

    \I__2165\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10137\
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__10143\,
            I => \config_register_latched_dec_inst.STATSRZ0Z_0\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__10140\,
            I => \config_register_latched_dec_inst.STATSRZ0Z_0\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__10137\,
            I => \config_register_latched_dec_inst.STATSRZ0Z_0\
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__10130\,
            I => \N__10127\
        );

    \I__2160\ : InMux
    port map (
            O => \N__10127\,
            I => \N__10124\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__10124\,
            I => \N__10120\
        );

    \I__2158\ : InMux
    port map (
            O => \N__10123\,
            I => \N__10117\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__10120\,
            I => \config_register_latched_dec_inst.STATCNF_1Z0Z_0\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__10117\,
            I => \config_register_latched_dec_inst.STATCNF_1Z0Z_0\
        );

    \I__2155\ : IoInMux
    port map (
            O => \N__10112\,
            I => \N__10109\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__10109\,
            I => \N__10106\
        );

    \I__2153\ : IoSpan4Mux
    port map (
            O => \N__10106\,
            I => \N__10102\
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__10105\,
            I => \N__10099\
        );

    \I__2151\ : Span4Mux_s2_h
    port map (
            O => \N__10102\,
            I => \N__10095\
        );

    \I__2150\ : InMux
    port map (
            O => \N__10099\,
            I => \N__10089\
        );

    \I__2149\ : InMux
    port map (
            O => \N__10098\,
            I => \N__10089\
        );

    \I__2148\ : Span4Mux_h
    port map (
            O => \N__10095\,
            I => \N__10075\
        );

    \I__2147\ : InMux
    port map (
            O => \N__10094\,
            I => \N__10064\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__10089\,
            I => \N__10061\
        );

    \I__2145\ : InMux
    port map (
            O => \N__10088\,
            I => \N__10050\
        );

    \I__2144\ : InMux
    port map (
            O => \N__10087\,
            I => \N__10050\
        );

    \I__2143\ : InMux
    port map (
            O => \N__10086\,
            I => \N__10050\
        );

    \I__2142\ : InMux
    port map (
            O => \N__10085\,
            I => \N__10050\
        );

    \I__2141\ : InMux
    port map (
            O => \N__10084\,
            I => \N__10050\
        );

    \I__2140\ : InMux
    port map (
            O => \N__10083\,
            I => \N__10047\
        );

    \I__2139\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10042\
        );

    \I__2138\ : InMux
    port map (
            O => \N__10081\,
            I => \N__10042\
        );

    \I__2137\ : InMux
    port map (
            O => \N__10080\,
            I => \N__10035\
        );

    \I__2136\ : InMux
    port map (
            O => \N__10079\,
            I => \N__10035\
        );

    \I__2135\ : InMux
    port map (
            O => \N__10078\,
            I => \N__10035\
        );

    \I__2134\ : Sp12to4
    port map (
            O => \N__10075\,
            I => \N__10032\
        );

    \I__2133\ : InMux
    port map (
            O => \N__10074\,
            I => \N__10021\
        );

    \I__2132\ : InMux
    port map (
            O => \N__10073\,
            I => \N__10021\
        );

    \I__2131\ : InMux
    port map (
            O => \N__10072\,
            I => \N__10021\
        );

    \I__2130\ : InMux
    port map (
            O => \N__10071\,
            I => \N__10021\
        );

    \I__2129\ : InMux
    port map (
            O => \N__10070\,
            I => \N__10021\
        );

    \I__2128\ : InMux
    port map (
            O => \N__10069\,
            I => \N__10014\
        );

    \I__2127\ : InMux
    port map (
            O => \N__10068\,
            I => \N__10014\
        );

    \I__2126\ : InMux
    port map (
            O => \N__10067\,
            I => \N__10014\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__10064\,
            I => \N__10011\
        );

    \I__2124\ : Span4Mux_v
    port map (
            O => \N__10061\,
            I => \N__10008\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__10050\,
            I => \N__9999\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__10047\,
            I => \N__9999\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__10042\,
            I => \N__9999\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__10035\,
            I => \N__9999\
        );

    \I__2119\ : Span12Mux_h
    port map (
            O => \N__10032\,
            I => \N__9996\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__10021\,
            I => \N__9991\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__10014\,
            I => \N__9991\
        );

    \I__2116\ : Span4Mux_v
    port map (
            O => \N__10011\,
            I => \N__9984\
        );

    \I__2115\ : Span4Mux_h
    port map (
            O => \N__10008\,
            I => \N__9984\
        );

    \I__2114\ : Span4Mux_v
    port map (
            O => \N__9999\,
            I => \N__9984\
        );

    \I__2113\ : Odrv12
    port map (
            O => \N__9996\,
            I => sel_output_c
        );

    \I__2112\ : Odrv12
    port map (
            O => \N__9991\,
            I => sel_output_c
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__9984\,
            I => sel_output_c
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__9977\,
            I => \N__9974\
        );

    \I__2109\ : InMux
    port map (
            O => \N__9974\,
            I => \N__9967\
        );

    \I__2108\ : InMux
    port map (
            O => \N__9973\,
            I => \N__9964\
        );

    \I__2107\ : InMux
    port map (
            O => \N__9972\,
            I => \N__9961\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9971\,
            I => \N__9956\
        );

    \I__2105\ : InMux
    port map (
            O => \N__9970\,
            I => \N__9956\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__9967\,
            I => \N__9951\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__9964\,
            I => \N__9951\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__9961\,
            I => \N__9948\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9956\,
            I => \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_2\
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__9951\,
            I => \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_2\
        );

    \I__2099\ : Odrv12
    port map (
            O => \N__9948\,
            I => \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_2\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9941\,
            I => \N__9937\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__9940\,
            I => \N__9933\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__9937\,
            I => \N__9928\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9936\,
            I => \N__9925\
        );

    \I__2094\ : InMux
    port map (
            O => \N__9933\,
            I => \N__9918\
        );

    \I__2093\ : InMux
    port map (
            O => \N__9932\,
            I => \N__9918\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9931\,
            I => \N__9918\
        );

    \I__2091\ : Odrv12
    port map (
            O => \N__9928\,
            I => \FSM_TEST_inst_RAPIDA.counter_dinZ1Z_1\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9925\,
            I => \FSM_TEST_inst_RAPIDA.counter_dinZ1Z_1\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__9918\,
            I => \FSM_TEST_inst_RAPIDA.counter_dinZ1Z_1\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__9911\,
            I => \N__9906\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__9910\,
            I => \N__9903\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__9909\,
            I => \N__9900\
        );

    \I__2085\ : InMux
    port map (
            O => \N__9906\,
            I => \N__9897\
        );

    \I__2084\ : InMux
    port map (
            O => \N__9903\,
            I => \N__9894\
        );

    \I__2083\ : InMux
    port map (
            O => \N__9900\,
            I => \N__9891\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__9897\,
            I => \N__9888\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__9894\,
            I => \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_3\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__9891\,
            I => \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_3\
        );

    \I__2079\ : Odrv12
    port map (
            O => \N__9888\,
            I => \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_3\
        );

    \I__2078\ : InMux
    port map (
            O => \N__9881\,
            I => \N__9874\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9880\,
            I => \N__9866\
        );

    \I__2076\ : InMux
    port map (
            O => \N__9879\,
            I => \N__9866\
        );

    \I__2075\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9866\
        );

    \I__2074\ : InMux
    port map (
            O => \N__9877\,
            I => \N__9863\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__9874\,
            I => \N__9860\
        );

    \I__2072\ : InMux
    port map (
            O => \N__9873\,
            I => \N__9857\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__9866\,
            I => \N__9854\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__9863\,
            I => \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_0\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__9860\,
            I => \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_0\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__9857\,
            I => \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_0\
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__9854\,
            I => \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_0\
        );

    \I__2066\ : InMux
    port map (
            O => \N__9845\,
            I => \N__9842\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9842\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_66\
        );

    \I__2064\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9836\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__9836\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_67\
        );

    \I__2062\ : InMux
    port map (
            O => \N__9833\,
            I => \N__9830\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__9830\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_45\
        );

    \I__2060\ : InMux
    port map (
            O => \N__9827\,
            I => \N__9824\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__9824\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_38\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9821\,
            I => \N__9818\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__9818\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_36\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9815\,
            I => \N__9812\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__9812\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_48\
        );

    \I__2054\ : InMux
    port map (
            O => \N__9809\,
            I => \N__9806\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9806\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_49\
        );

    \I__2052\ : InMux
    port map (
            O => \N__9803\,
            I => \N__9800\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__9800\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_33\
        );

    \I__2050\ : InMux
    port map (
            O => \N__9797\,
            I => \N__9794\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9794\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_34\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9791\,
            I => \N__9788\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__9788\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_10\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9785\,
            I => \N__9782\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__9782\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_74\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9779\,
            I => \N__9776\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__9776\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_13\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9773\,
            I => \N__9770\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__9770\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_14\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9767\,
            I => \N__9764\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__9764\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_15\
        );

    \I__2038\ : InMux
    port map (
            O => \N__9761\,
            I => \N__9758\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__9758\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_16\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9752\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__9752\,
            I => \N__9749\
        );

    \I__2034\ : Odrv4
    port map (
            O => \N__9749\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_17\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9746\,
            I => \N__9743\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__9743\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_65\
        );

    \I__2031\ : InMux
    port map (
            O => \N__9740\,
            I => \N__9737\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9737\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_35\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9734\,
            I => \N__9731\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__9731\,
            I => \N__9728\
        );

    \I__2027\ : Odrv4
    port map (
            O => \N__9728\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_80\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9725\,
            I => \N__9722\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__9722\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_81\
        );

    \I__2024\ : InMux
    port map (
            O => \N__9719\,
            I => \N__9716\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__9716\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_32\
        );

    \I__2022\ : InMux
    port map (
            O => \N__9713\,
            I => \N__9710\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9710\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_39\
        );

    \I__2020\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9704\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__9704\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_46\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9701\,
            I => \N__9698\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__9698\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_47\
        );

    \I__2016\ : InMux
    port map (
            O => \N__9695\,
            I => \N__9692\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__9692\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_40\
        );

    \I__2014\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9686\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__9686\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_55\
        );

    \I__2012\ : InMux
    port map (
            O => \N__9683\,
            I => \N__9680\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__9680\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_56\
        );

    \I__2010\ : InMux
    port map (
            O => \N__9677\,
            I => \N__9674\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__9674\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_83\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__9671\,
            I => \N__9668\
        );

    \I__2007\ : InMux
    port map (
            O => \N__9668\,
            I => \N__9665\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__9665\,
            I => \N__9662\
        );

    \I__2005\ : Span4Mux_h
    port map (
            O => \N__9662\,
            I => \N__9659\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__9659\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_87\
        );

    \I__2003\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9653\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__9653\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_84\
        );

    \I__2001\ : InMux
    port map (
            O => \N__9650\,
            I => \N__9647\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9647\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_85\
        );

    \I__1999\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9641\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__9641\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_86\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9638\,
            I => \N__9635\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__9635\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_82\
        );

    \I__1995\ : InMux
    port map (
            O => \N__9632\,
            I => \N__9629\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__9629\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_29\
        );

    \I__1993\ : InMux
    port map (
            O => \N__9626\,
            I => \N__9623\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__9623\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_30\
        );

    \I__1991\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9617\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__9617\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_75\
        );

    \I__1989\ : InMux
    port map (
            O => \N__9614\,
            I => \N__9611\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__9611\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_60\
        );

    \I__1987\ : InMux
    port map (
            O => \N__9608\,
            I => \N__9605\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__9605\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_58\
        );

    \I__1985\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9599\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__9599\,
            I => \N__9596\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__9596\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_7\
        );

    \I__1982\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9590\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__9590\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_8\
        );

    \I__1980\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9584\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__9584\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_9\
        );

    \I__1978\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9578\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__9578\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_57\
        );

    \I__1976\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9572\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__9572\,
            I => \N__9569\
        );

    \I__1974\ : Span4Mux_h
    port map (
            O => \N__9569\,
            I => \N__9566\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__9566\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_79\
        );

    \I__1972\ : InMux
    port map (
            O => \N__9563\,
            I => \N__9557\
        );

    \I__1971\ : InMux
    port map (
            O => \N__9562\,
            I => \N__9557\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__9557\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_7\
        );

    \I__1969\ : InMux
    port map (
            O => \N__9554\,
            I => \N__9548\
        );

    \I__1968\ : InMux
    port map (
            O => \N__9553\,
            I => \N__9548\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__9548\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_5\
        );

    \I__1966\ : InMux
    port map (
            O => \N__9545\,
            I => \N__9539\
        );

    \I__1965\ : InMux
    port map (
            O => \N__9544\,
            I => \N__9539\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__9539\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_6\
        );

    \I__1963\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9532\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9535\,
            I => \N__9529\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__9532\,
            I => \N__9522\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__9529\,
            I => \N__9522\
        );

    \I__1959\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9517\
        );

    \I__1958\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9517\
        );

    \I__1957\ : Span4Mux_h
    port map (
            O => \N__9522\,
            I => \N__9514\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__9517\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_8\
        );

    \I__1955\ : Odrv4
    port map (
            O => \N__9514\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_8\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__9509\,
            I => \N__9506\
        );

    \I__1953\ : InMux
    port map (
            O => \N__9506\,
            I => \N__9500\
        );

    \I__1952\ : InMux
    port map (
            O => \N__9505\,
            I => \N__9500\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__9500\,
            I => \N__9495\
        );

    \I__1950\ : InMux
    port map (
            O => \N__9499\,
            I => \N__9492\
        );

    \I__1949\ : InMux
    port map (
            O => \N__9498\,
            I => \N__9489\
        );

    \I__1948\ : Span4Mux_h
    port map (
            O => \N__9495\,
            I => \N__9486\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__9492\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_9\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__9489\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_9\
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__9486\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_9\
        );

    \I__1944\ : CEMux
    port map (
            O => \N__9479\,
            I => \N__9475\
        );

    \I__1943\ : CEMux
    port map (
            O => \N__9478\,
            I => \N__9472\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__9475\,
            I => \N__9469\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__9472\,
            I => \N__9466\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__9469\,
            I => \N__9463\
        );

    \I__1939\ : Span4Mux_v
    port map (
            O => \N__9466\,
            I => \N__9460\
        );

    \I__1938\ : Odrv4
    port map (
            O => \N__9463\,
            I => \flag_output_0_ret_RNI1E8NZ0Z2\
        );

    \I__1937\ : Odrv4
    port map (
            O => \N__9460\,
            I => \flag_output_0_ret_RNI1E8NZ0Z2\
        );

    \I__1936\ : InMux
    port map (
            O => \N__9455\,
            I => \N__9452\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__9452\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_51\
        );

    \I__1934\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__9446\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_52\
        );

    \I__1932\ : InMux
    port map (
            O => \N__9443\,
            I => \N__9440\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__9440\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_53\
        );

    \I__1930\ : InMux
    port map (
            O => \N__9437\,
            I => \N__9434\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__9434\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_31\
        );

    \I__1928\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__9428\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_50\
        );

    \I__1926\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9421\
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__9424\,
            I => \N__9415\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__9421\,
            I => \N__9408\
        );

    \I__1923\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9405\
        );

    \I__1922\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9394\
        );

    \I__1921\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9394\
        );

    \I__1920\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9394\
        );

    \I__1919\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9394\
        );

    \I__1918\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9394\
        );

    \I__1917\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9391\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__9411\,
            I => \N__9388\
        );

    \I__1915\ : Span4Mux_h
    port map (
            O => \N__9408\,
            I => \N__9382\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__9405\,
            I => \N__9382\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__9394\,
            I => \N__9377\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__9391\,
            I => \N__9377\
        );

    \I__1911\ : InMux
    port map (
            O => \N__9388\,
            I => \N__9374\
        );

    \I__1910\ : InMux
    port map (
            O => \N__9387\,
            I => \N__9371\
        );

    \I__1909\ : Span4Mux_v
    port map (
            O => \N__9382\,
            I => \N__9368\
        );

    \I__1908\ : Span4Mux_h
    port map (
            O => \N__9377\,
            I => \N__9365\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__9374\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fastZ0Z_1\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__9371\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fastZ0Z_1\
        );

    \I__1905\ : Odrv4
    port map (
            O => \N__9368\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fastZ0Z_1\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__9365\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fastZ0Z_1\
        );

    \I__1903\ : InMux
    port map (
            O => \N__9356\,
            I => \N__9353\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__9353\,
            I => \N__9350\
        );

    \I__1901\ : Odrv12
    port map (
            O => \N__9350\,
            I => \FSM_TEST_inst_slow.CLK_uC_6kZ0Z_0\
        );

    \I__1900\ : InMux
    port map (
            O => \N__9347\,
            I => \N__9344\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__9344\,
            I => \N__9340\
        );

    \I__1898\ : InMux
    port map (
            O => \N__9343\,
            I => \N__9337\
        );

    \I__1897\ : Odrv4
    port map (
            O => \N__9340\,
            I => \CLK_uC_6l_0\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__9337\,
            I => \CLK_uC_6l_0\
        );

    \I__1895\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9326\
        );

    \I__1894\ : InMux
    port map (
            O => \N__9331\,
            I => \N__9326\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__9326\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_3\
        );

    \I__1892\ : InMux
    port map (
            O => \N__9323\,
            I => \N__9317\
        );

    \I__1891\ : InMux
    port map (
            O => \N__9322\,
            I => \N__9317\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__9317\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_4\
        );

    \I__1889\ : InMux
    port map (
            O => \N__9314\,
            I => \N__9310\
        );

    \I__1888\ : InMux
    port map (
            O => \N__9313\,
            I => \N__9307\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__9310\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_1\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__9307\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_1\
        );

    \I__1885\ : InMux
    port map (
            O => \N__9302\,
            I => \N__9296\
        );

    \I__1884\ : InMux
    port map (
            O => \N__9301\,
            I => \N__9296\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__9296\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_2\
        );

    \I__1882\ : InMux
    port map (
            O => \N__9293\,
            I => \N__9284\
        );

    \I__1881\ : InMux
    port map (
            O => \N__9292\,
            I => \N__9281\
        );

    \I__1880\ : InMux
    port map (
            O => \N__9291\,
            I => \N__9270\
        );

    \I__1879\ : InMux
    port map (
            O => \N__9290\,
            I => \N__9270\
        );

    \I__1878\ : InMux
    port map (
            O => \N__9289\,
            I => \N__9270\
        );

    \I__1877\ : InMux
    port map (
            O => \N__9288\,
            I => \N__9270\
        );

    \I__1876\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9270\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__9284\,
            I => \N__9265\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__9281\,
            I => \N__9265\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__9270\,
            I => \FSM_TEST_inst_slow.current_state_RNI9C3K2Z0Z_1\
        );

    \I__1872\ : Odrv12
    port map (
            O => \N__9265\,
            I => \FSM_TEST_inst_slow.current_state_RNI9C3K2Z0Z_1\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__9260\,
            I => \N__9256\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__9259\,
            I => \N__9251\
        );

    \I__1869\ : InMux
    port map (
            O => \N__9256\,
            I => \N__9247\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__9255\,
            I => \N__9244\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__9254\,
            I => \N__9241\
        );

    \I__1866\ : InMux
    port map (
            O => \N__9251\,
            I => \N__9236\
        );

    \I__1865\ : InMux
    port map (
            O => \N__9250\,
            I => \N__9233\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__9247\,
            I => \N__9230\
        );

    \I__1863\ : InMux
    port map (
            O => \N__9244\,
            I => \N__9221\
        );

    \I__1862\ : InMux
    port map (
            O => \N__9241\,
            I => \N__9221\
        );

    \I__1861\ : InMux
    port map (
            O => \N__9240\,
            I => \N__9221\
        );

    \I__1860\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9221\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__9236\,
            I => \N__9216\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__9233\,
            I => \N__9216\
        );

    \I__1857\ : Span4Mux_h
    port map (
            O => \N__9230\,
            I => \N__9213\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__9221\,
            I => \FSM_TEST_inst_slow.current_state_d_i_2\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__9216\,
            I => \FSM_TEST_inst_slow.current_state_d_i_2\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__9213\,
            I => \FSM_TEST_inst_slow.current_state_d_i_2\
        );

    \I__1853\ : InMux
    port map (
            O => \N__9206\,
            I => \N__9203\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__9203\,
            I => \N__9200\
        );

    \I__1851\ : Odrv4
    port map (
            O => \N__9200\,
            I => \FSM_TEST_inst_slow.counter_stat_cry_4_THRU_CO\
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__9197\,
            I => \N__9193\
        );

    \I__1849\ : InMux
    port map (
            O => \N__9196\,
            I => \N__9189\
        );

    \I__1848\ : InMux
    port map (
            O => \N__9193\,
            I => \N__9186\
        );

    \I__1847\ : InMux
    port map (
            O => \N__9192\,
            I => \N__9183\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__9189\,
            I => \N__9175\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__9186\,
            I => \N__9175\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__9183\,
            I => \N__9175\
        );

    \I__1843\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9172\
        );

    \I__1842\ : Span4Mux_h
    port map (
            O => \N__9175\,
            I => \N__9169\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__9172\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_5\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__9169\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_5\
        );

    \I__1839\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9153\
        );

    \I__1838\ : InMux
    port map (
            O => \N__9163\,
            I => \N__9153\
        );

    \I__1837\ : InMux
    port map (
            O => \N__9162\,
            I => \N__9153\
        );

    \I__1836\ : InMux
    port map (
            O => \N__9161\,
            I => \N__9148\
        );

    \I__1835\ : InMux
    port map (
            O => \N__9160\,
            I => \N__9148\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__9153\,
            I => \N__9145\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__9148\,
            I => \divisor_inst_2.counterZ0Z_1\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__9145\,
            I => \divisor_inst_2.counterZ0Z_1\
        );

    \I__1831\ : CascadeMux
    port map (
            O => \N__9140\,
            I => \N__9136\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__9139\,
            I => \N__9131\
        );

    \I__1829\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9122\
        );

    \I__1828\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9122\
        );

    \I__1827\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9122\
        );

    \I__1826\ : InMux
    port map (
            O => \N__9131\,
            I => \N__9115\
        );

    \I__1825\ : InMux
    port map (
            O => \N__9130\,
            I => \N__9115\
        );

    \I__1824\ : InMux
    port map (
            O => \N__9129\,
            I => \N__9115\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__9122\,
            I => \divisor_inst_2.counterZ0Z_0\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__9115\,
            I => \divisor_inst_2.counterZ0Z_0\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__9110\,
            I => \N__9104\
        );

    \I__1820\ : CascadeMux
    port map (
            O => \N__9109\,
            I => \N__9101\
        );

    \I__1819\ : InMux
    port map (
            O => \N__9108\,
            I => \N__9098\
        );

    \I__1818\ : InMux
    port map (
            O => \N__9107\,
            I => \N__9091\
        );

    \I__1817\ : InMux
    port map (
            O => \N__9104\,
            I => \N__9091\
        );

    \I__1816\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9091\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__9098\,
            I => \divisor_inst_2.counterZ0Z_2\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__9091\,
            I => \divisor_inst_2.counterZ0Z_2\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__9086\,
            I => \N__9082\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__9085\,
            I => \N__9078\
        );

    \I__1811\ : InMux
    port map (
            O => \N__9082\,
            I => \N__9075\
        );

    \I__1810\ : InMux
    port map (
            O => \N__9081\,
            I => \N__9072\
        );

    \I__1809\ : InMux
    port map (
            O => \N__9078\,
            I => \N__9069\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__9075\,
            I => \FSM_TEST_inst_RAPIDA.aux_selection_fast_0\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__9072\,
            I => \FSM_TEST_inst_RAPIDA.aux_selection_fast_0\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__9069\,
            I => \FSM_TEST_inst_RAPIDA.aux_selection_fast_0\
        );

    \I__1805\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9057\
        );

    \I__1804\ : InMux
    port map (
            O => \N__9061\,
            I => \N__9052\
        );

    \I__1803\ : InMux
    port map (
            O => \N__9060\,
            I => \N__9052\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__9057\,
            I => \N__9038\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__9052\,
            I => \N__9035\
        );

    \I__1800\ : InMux
    port map (
            O => \N__9051\,
            I => \N__9030\
        );

    \I__1799\ : InMux
    port map (
            O => \N__9050\,
            I => \N__9030\
        );

    \I__1798\ : InMux
    port map (
            O => \N__9049\,
            I => \N__8995\
        );

    \I__1797\ : InMux
    port map (
            O => \N__9048\,
            I => \N__8995\
        );

    \I__1796\ : InMux
    port map (
            O => \N__9047\,
            I => \N__8995\
        );

    \I__1795\ : InMux
    port map (
            O => \N__9046\,
            I => \N__8992\
        );

    \I__1794\ : InMux
    port map (
            O => \N__9045\,
            I => \N__8989\
        );

    \I__1793\ : InMux
    port map (
            O => \N__9044\,
            I => \N__8947\
        );

    \I__1792\ : InMux
    port map (
            O => \N__9043\,
            I => \N__8942\
        );

    \I__1791\ : InMux
    port map (
            O => \N__9042\,
            I => \N__8942\
        );

    \I__1790\ : InMux
    port map (
            O => \N__9041\,
            I => \N__8927\
        );

    \I__1789\ : Span4Mux_v
    port map (
            O => \N__9038\,
            I => \N__8920\
        );

    \I__1788\ : Span4Mux_h
    port map (
            O => \N__9035\,
            I => \N__8920\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__9030\,
            I => \N__8920\
        );

    \I__1786\ : InMux
    port map (
            O => \N__9029\,
            I => \N__8909\
        );

    \I__1785\ : InMux
    port map (
            O => \N__9028\,
            I => \N__8909\
        );

    \I__1784\ : InMux
    port map (
            O => \N__9027\,
            I => \N__8909\
        );

    \I__1783\ : InMux
    port map (
            O => \N__9026\,
            I => \N__8909\
        );

    \I__1782\ : InMux
    port map (
            O => \N__9025\,
            I => \N__8909\
        );

    \I__1781\ : InMux
    port map (
            O => \N__9024\,
            I => \N__8898\
        );

    \I__1780\ : InMux
    port map (
            O => \N__9023\,
            I => \N__8898\
        );

    \I__1779\ : InMux
    port map (
            O => \N__9022\,
            I => \N__8898\
        );

    \I__1778\ : InMux
    port map (
            O => \N__9021\,
            I => \N__8898\
        );

    \I__1777\ : InMux
    port map (
            O => \N__9020\,
            I => \N__8898\
        );

    \I__1776\ : InMux
    port map (
            O => \N__9019\,
            I => \N__8883\
        );

    \I__1775\ : InMux
    port map (
            O => \N__9018\,
            I => \N__8883\
        );

    \I__1774\ : InMux
    port map (
            O => \N__9017\,
            I => \N__8883\
        );

    \I__1773\ : InMux
    port map (
            O => \N__9016\,
            I => \N__8883\
        );

    \I__1772\ : InMux
    port map (
            O => \N__9015\,
            I => \N__8883\
        );

    \I__1771\ : InMux
    port map (
            O => \N__9014\,
            I => \N__8883\
        );

    \I__1770\ : InMux
    port map (
            O => \N__9013\,
            I => \N__8883\
        );

    \I__1769\ : InMux
    port map (
            O => \N__9012\,
            I => \N__8880\
        );

    \I__1768\ : InMux
    port map (
            O => \N__9011\,
            I => \N__8863\
        );

    \I__1767\ : InMux
    port map (
            O => \N__9010\,
            I => \N__8863\
        );

    \I__1766\ : InMux
    port map (
            O => \N__9009\,
            I => \N__8863\
        );

    \I__1765\ : InMux
    port map (
            O => \N__9008\,
            I => \N__8863\
        );

    \I__1764\ : InMux
    port map (
            O => \N__9007\,
            I => \N__8863\
        );

    \I__1763\ : InMux
    port map (
            O => \N__9006\,
            I => \N__8863\
        );

    \I__1762\ : InMux
    port map (
            O => \N__9005\,
            I => \N__8863\
        );

    \I__1761\ : InMux
    port map (
            O => \N__9004\,
            I => \N__8863\
        );

    \I__1760\ : InMux
    port map (
            O => \N__9003\,
            I => \N__8858\
        );

    \I__1759\ : InMux
    port map (
            O => \N__9002\,
            I => \N__8858\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__8995\,
            I => \N__8851\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__8992\,
            I => \N__8848\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8989\,
            I => \N__8845\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8988\,
            I => \N__8834\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8987\,
            I => \N__8834\
        );

    \I__1753\ : InMux
    port map (
            O => \N__8986\,
            I => \N__8834\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8985\,
            I => \N__8834\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8834\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8983\,
            I => \N__8827\
        );

    \I__1749\ : InMux
    port map (
            O => \N__8982\,
            I => \N__8827\
        );

    \I__1748\ : InMux
    port map (
            O => \N__8981\,
            I => \N__8827\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8980\,
            I => \N__8824\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8979\,
            I => \N__8817\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8978\,
            I => \N__8817\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8817\
        );

    \I__1743\ : InMux
    port map (
            O => \N__8976\,
            I => \N__8804\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8804\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8974\,
            I => \N__8804\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8973\,
            I => \N__8804\
        );

    \I__1739\ : InMux
    port map (
            O => \N__8972\,
            I => \N__8804\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8971\,
            I => \N__8804\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8789\
        );

    \I__1736\ : InMux
    port map (
            O => \N__8969\,
            I => \N__8789\
        );

    \I__1735\ : InMux
    port map (
            O => \N__8968\,
            I => \N__8789\
        );

    \I__1734\ : InMux
    port map (
            O => \N__8967\,
            I => \N__8789\
        );

    \I__1733\ : InMux
    port map (
            O => \N__8966\,
            I => \N__8789\
        );

    \I__1732\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8789\
        );

    \I__1731\ : InMux
    port map (
            O => \N__8964\,
            I => \N__8789\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8963\,
            I => \N__8778\
        );

    \I__1729\ : InMux
    port map (
            O => \N__8962\,
            I => \N__8778\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8961\,
            I => \N__8778\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8960\,
            I => \N__8778\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8959\,
            I => \N__8778\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8958\,
            I => \N__8769\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8957\,
            I => \N__8769\
        );

    \I__1723\ : InMux
    port map (
            O => \N__8956\,
            I => \N__8769\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8955\,
            I => \N__8769\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8954\,
            I => \N__8765\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8953\,
            I => \N__8756\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8952\,
            I => \N__8756\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8951\,
            I => \N__8756\
        );

    \I__1717\ : InMux
    port map (
            O => \N__8950\,
            I => \N__8756\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__8947\,
            I => \N__8751\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8942\,
            I => \N__8751\
        );

    \I__1714\ : InMux
    port map (
            O => \N__8941\,
            I => \N__8742\
        );

    \I__1713\ : InMux
    port map (
            O => \N__8940\,
            I => \N__8742\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8939\,
            I => \N__8742\
        );

    \I__1711\ : InMux
    port map (
            O => \N__8938\,
            I => \N__8742\
        );

    \I__1710\ : InMux
    port map (
            O => \N__8937\,
            I => \N__8725\
        );

    \I__1709\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8725\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8935\,
            I => \N__8725\
        );

    \I__1707\ : InMux
    port map (
            O => \N__8934\,
            I => \N__8725\
        );

    \I__1706\ : InMux
    port map (
            O => \N__8933\,
            I => \N__8725\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8932\,
            I => \N__8725\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8931\,
            I => \N__8725\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8930\,
            I => \N__8725\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__8927\,
            I => \N__8698\
        );

    \I__1701\ : Span4Mux_h
    port map (
            O => \N__8920\,
            I => \N__8698\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8909\,
            I => \N__8698\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__8898\,
            I => \N__8698\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__8883\,
            I => \N__8698\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__8880\,
            I => \N__8695\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__8863\,
            I => \N__8690\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8858\,
            I => \N__8690\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8857\,
            I => \N__8681\
        );

    \I__1693\ : InMux
    port map (
            O => \N__8856\,
            I => \N__8681\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8855\,
            I => \N__8681\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8854\,
            I => \N__8681\
        );

    \I__1690\ : Span4Mux_v
    port map (
            O => \N__8851\,
            I => \N__8670\
        );

    \I__1689\ : Span4Mux_h
    port map (
            O => \N__8848\,
            I => \N__8670\
        );

    \I__1688\ : Span4Mux_v
    port map (
            O => \N__8845\,
            I => \N__8670\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__8834\,
            I => \N__8670\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__8827\,
            I => \N__8670\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__8824\,
            I => \N__8657\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__8817\,
            I => \N__8657\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8804\,
            I => \N__8657\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__8789\,
            I => \N__8657\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__8778\,
            I => \N__8657\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__8769\,
            I => \N__8657\
        );

    \I__1679\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8654\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__8765\,
            I => \N__8645\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__8756\,
            I => \N__8645\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__8751\,
            I => \N__8640\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__8742\,
            I => \N__8640\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8725\,
            I => \N__8637\
        );

    \I__1673\ : InMux
    port map (
            O => \N__8724\,
            I => \N__8626\
        );

    \I__1672\ : InMux
    port map (
            O => \N__8723\,
            I => \N__8626\
        );

    \I__1671\ : InMux
    port map (
            O => \N__8722\,
            I => \N__8626\
        );

    \I__1670\ : InMux
    port map (
            O => \N__8721\,
            I => \N__8626\
        );

    \I__1669\ : InMux
    port map (
            O => \N__8720\,
            I => \N__8626\
        );

    \I__1668\ : InMux
    port map (
            O => \N__8719\,
            I => \N__8611\
        );

    \I__1667\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8611\
        );

    \I__1666\ : InMux
    port map (
            O => \N__8717\,
            I => \N__8611\
        );

    \I__1665\ : InMux
    port map (
            O => \N__8716\,
            I => \N__8611\
        );

    \I__1664\ : InMux
    port map (
            O => \N__8715\,
            I => \N__8611\
        );

    \I__1663\ : InMux
    port map (
            O => \N__8714\,
            I => \N__8611\
        );

    \I__1662\ : InMux
    port map (
            O => \N__8713\,
            I => \N__8611\
        );

    \I__1661\ : InMux
    port map (
            O => \N__8712\,
            I => \N__8604\
        );

    \I__1660\ : InMux
    port map (
            O => \N__8711\,
            I => \N__8604\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8710\,
            I => \N__8604\
        );

    \I__1658\ : InMux
    port map (
            O => \N__8709\,
            I => \N__8601\
        );

    \I__1657\ : Span4Mux_v
    port map (
            O => \N__8698\,
            I => \N__8592\
        );

    \I__1656\ : Span4Mux_v
    port map (
            O => \N__8695\,
            I => \N__8592\
        );

    \I__1655\ : Span4Mux_v
    port map (
            O => \N__8690\,
            I => \N__8592\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__8681\,
            I => \N__8592\
        );

    \I__1653\ : Span4Mux_h
    port map (
            O => \N__8670\,
            I => \N__8585\
        );

    \I__1652\ : Span4Mux_v
    port map (
            O => \N__8657\,
            I => \N__8585\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__8654\,
            I => \N__8585\
        );

    \I__1650\ : InMux
    port map (
            O => \N__8653\,
            I => \N__8576\
        );

    \I__1649\ : InMux
    port map (
            O => \N__8652\,
            I => \N__8576\
        );

    \I__1648\ : InMux
    port map (
            O => \N__8651\,
            I => \N__8576\
        );

    \I__1647\ : InMux
    port map (
            O => \N__8650\,
            I => \N__8576\
        );

    \I__1646\ : Odrv12
    port map (
            O => \N__8645\,
            I => \FSM_TEST_inst_slow.current_stateZ1Z_0\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__8640\,
            I => \FSM_TEST_inst_slow.current_stateZ1Z_0\
        );

    \I__1644\ : Odrv4
    port map (
            O => \N__8637\,
            I => \FSM_TEST_inst_slow.current_stateZ1Z_0\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__8626\,
            I => \FSM_TEST_inst_slow.current_stateZ1Z_0\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__8611\,
            I => \FSM_TEST_inst_slow.current_stateZ1Z_0\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__8604\,
            I => \FSM_TEST_inst_slow.current_stateZ1Z_0\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__8601\,
            I => \FSM_TEST_inst_slow.current_stateZ1Z_0\
        );

    \I__1639\ : Odrv4
    port map (
            O => \N__8592\,
            I => \FSM_TEST_inst_slow.current_stateZ1Z_0\
        );

    \I__1638\ : Odrv4
    port map (
            O => \N__8585\,
            I => \FSM_TEST_inst_slow.current_stateZ1Z_0\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__8576\,
            I => \FSM_TEST_inst_slow.current_stateZ1Z_0\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__8555\,
            I => \N__8552\
        );

    \I__1635\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8549\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__8549\,
            I => \counter_RNIFD27_2\
        );

    \I__1633\ : InMux
    port map (
            O => \N__8546\,
            I => \N__8543\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__8543\,
            I => \N__8540\
        );

    \I__1631\ : Span4Mux_h
    port map (
            O => \N__8540\,
            I => \N__8537\
        );

    \I__1630\ : Span4Mux_h
    port map (
            O => \N__8537\,
            I => \N__8530\
        );

    \I__1629\ : InMux
    port map (
            O => \N__8536\,
            I => \N__8527\
        );

    \I__1628\ : InMux
    port map (
            O => \N__8535\,
            I => \N__8520\
        );

    \I__1627\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8520\
        );

    \I__1626\ : InMux
    port map (
            O => \N__8533\,
            I => \N__8520\
        );

    \I__1625\ : Odrv4
    port map (
            O => \N__8530\,
            I => clk_continuous_slow
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__8527\,
            I => clk_continuous_slow
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__8520\,
            I => clk_continuous_slow
        );

    \I__1622\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8509\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8506\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__8509\,
            I => \N__8503\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__8506\,
            I => \FSM_TEST_inst_slow.aux_selection_slow_0\
        );

    \I__1618\ : Odrv4
    port map (
            O => \N__8503\,
            I => \FSM_TEST_inst_slow.aux_selection_slow_0\
        );

    \I__1617\ : CascadeMux
    port map (
            O => \N__8498\,
            I => \N__8493\
        );

    \I__1616\ : InMux
    port map (
            O => \N__8497\,
            I => \N__8490\
        );

    \I__1615\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8487\
        );

    \I__1614\ : InMux
    port map (
            O => \N__8493\,
            I => \N__8483\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__8490\,
            I => \N__8478\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__8487\,
            I => \N__8478\
        );

    \I__1611\ : InMux
    port map (
            O => \N__8486\,
            I => \N__8475\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__8483\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_fastZ0Z_1\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__8478\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_fastZ0Z_1\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__8475\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_fastZ0Z_1\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__8468\,
            I => \N__8464\
        );

    \I__1606\ : InMux
    port map (
            O => \N__8467\,
            I => \N__8457\
        );

    \I__1605\ : InMux
    port map (
            O => \N__8464\,
            I => \N__8457\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__8463\,
            I => \N__8451\
        );

    \I__1603\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8447\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__8457\,
            I => \N__8444\
        );

    \I__1601\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8441\
        );

    \I__1600\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8434\
        );

    \I__1599\ : InMux
    port map (
            O => \N__8454\,
            I => \N__8434\
        );

    \I__1598\ : InMux
    port map (
            O => \N__8451\,
            I => \N__8434\
        );

    \I__1597\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8429\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__8447\,
            I => \N__8420\
        );

    \I__1595\ : Span4Mux_v
    port map (
            O => \N__8444\,
            I => \N__8420\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__8441\,
            I => \N__8420\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__8434\,
            I => \N__8420\
        );

    \I__1592\ : InMux
    port map (
            O => \N__8433\,
            I => \N__8415\
        );

    \I__1591\ : InMux
    port map (
            O => \N__8432\,
            I => \N__8415\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__8429\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_1_repZ0Z1\
        );

    \I__1589\ : Odrv4
    port map (
            O => \N__8420\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_1_repZ0Z1\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__8415\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_1_repZ0Z1\
        );

    \I__1587\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8405\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__8405\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_76\
        );

    \I__1585\ : InMux
    port map (
            O => \N__8402\,
            I => \N__8399\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__8399\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_54\
        );

    \I__1583\ : InMux
    port map (
            O => \N__8396\,
            I => \N__8393\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__8393\,
            I => \FSM_TEST_inst_RAPIDA.CLK_uC_2Z0Z_0\
        );

    \I__1581\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8387\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__8387\,
            I => \FSM_TEST_inst_RAPIDA.CLK_uC_6bZ0Z_0\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__8384\,
            I => \N__8380\
        );

    \I__1578\ : InMux
    port map (
            O => \N__8383\,
            I => \N__8375\
        );

    \I__1577\ : InMux
    port map (
            O => \N__8380\,
            I => \N__8375\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__8375\,
            I => \FSM_TEST_inst_RAPIDA.CLK_uCZ0\
        );

    \I__1575\ : InMux
    port map (
            O => \N__8372\,
            I => \N__8369\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__8369\,
            I => \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5DZ0Z1\
        );

    \I__1573\ : InMux
    port map (
            O => \N__8366\,
            I => \N__8362\
        );

    \I__1572\ : InMux
    port map (
            O => \N__8365\,
            I => \N__8359\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__8362\,
            I => \N_3_0\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__8359\,
            I => \N_3_0\
        );

    \I__1569\ : InMux
    port map (
            O => \N__8354\,
            I => \N__8345\
        );

    \I__1568\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8345\
        );

    \I__1567\ : InMux
    port map (
            O => \N__8352\,
            I => \N__8342\
        );

    \I__1566\ : InMux
    port map (
            O => \N__8351\,
            I => \N__8339\
        );

    \I__1565\ : InMux
    port map (
            O => \N__8350\,
            I => \N__8336\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__8345\,
            I => \N_4_0\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__8342\,
            I => \N_4_0\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__8339\,
            I => \N_4_0\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__8336\,
            I => \N_4_0\
        );

    \I__1560\ : InMux
    port map (
            O => \N__8327\,
            I => \N__8323\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__8326\,
            I => \N__8320\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__8323\,
            I => \N__8317\
        );

    \I__1557\ : InMux
    port map (
            O => \N__8320\,
            I => \N__8314\
        );

    \I__1556\ : Span4Mux_v
    port map (
            O => \N__8317\,
            I => \N__8309\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__8314\,
            I => \N__8309\
        );

    \I__1554\ : Span4Mux_h
    port map (
            O => \N__8309\,
            I => \N__8306\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__8306\,
            I => \CLK_uC_6c_0\
        );

    \I__1552\ : IoInMux
    port map (
            O => \N__8303\,
            I => \N__8300\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__8300\,
            I => \N__8297\
        );

    \I__1550\ : Span4Mux_s1_v
    port map (
            O => \N__8297\,
            I => \N__8294\
        );

    \I__1549\ : Span4Mux_v
    port map (
            O => \N__8294\,
            I => \N__8291\
        );

    \I__1548\ : Sp12to4
    port map (
            O => \N__8291\,
            I => \N__8287\
        );

    \I__1547\ : InMux
    port map (
            O => \N__8290\,
            I => \N__8284\
        );

    \I__1546\ : Span12Mux_h
    port map (
            O => \N__8287\,
            I => \N__8281\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__8284\,
            I => \N__8278\
        );

    \I__1544\ : Odrv12
    port map (
            O => \N__8281\,
            I => clk_output_c
        );

    \I__1543\ : Odrv4
    port map (
            O => \N__8278\,
            I => clk_output_c
        );

    \I__1542\ : InMux
    port map (
            O => \N__8273\,
            I => \N__8270\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__8270\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_6\
        );

    \I__1540\ : InMux
    port map (
            O => \N__8267\,
            I => \N__8264\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__8264\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_7\
        );

    \I__1538\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8258\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__8258\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_8\
        );

    \I__1536\ : InMux
    port map (
            O => \N__8255\,
            I => \N__8252\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__8252\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_9\
        );

    \I__1534\ : InMux
    port map (
            O => \N__8249\,
            I => \N__8246\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__8246\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_11\
        );

    \I__1532\ : InMux
    port map (
            O => \N__8243\,
            I => \N__8240\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__8240\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_12\
        );

    \I__1530\ : CEMux
    port map (
            O => \N__8237\,
            I => \N__8234\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__8234\,
            I => \N__8229\
        );

    \I__1528\ : CEMux
    port map (
            O => \N__8233\,
            I => \N__8226\
        );

    \I__1527\ : CEMux
    port map (
            O => \N__8232\,
            I => \N__8223\
        );

    \I__1526\ : Span4Mux_h
    port map (
            O => \N__8229\,
            I => \N__8218\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__8226\,
            I => \N__8218\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__8223\,
            I => \N__8215\
        );

    \I__1523\ : Odrv4
    port map (
            O => \N__8218\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_RNI78E11Z0Z_1\
        );

    \I__1522\ : Odrv12
    port map (
            O => \N__8215\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_RNI78E11Z0Z_1\
        );

    \I__1521\ : InMux
    port map (
            O => \N__8210\,
            I => \N__8207\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__8207\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_27\
        );

    \I__1519\ : InMux
    port map (
            O => \N__8204\,
            I => \N__8201\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__8201\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_28\
        );

    \I__1517\ : InMux
    port map (
            O => \N__8198\,
            I => \N__8195\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__8195\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_59\
        );

    \I__1515\ : InMux
    port map (
            O => \N__8192\,
            I => \N__8186\
        );

    \I__1514\ : InMux
    port map (
            O => \N__8191\,
            I => \N__8186\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__8186\,
            I => \N__8183\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__8183\,
            I => \FSM_TEST_inst_RAPIDA.N_101_0\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__8180\,
            I => \N__8176\
        );

    \I__1510\ : InMux
    port map (
            O => \N__8179\,
            I => \N__8172\
        );

    \I__1509\ : InMux
    port map (
            O => \N__8176\,
            I => \N__8169\
        );

    \I__1508\ : InMux
    port map (
            O => \N__8175\,
            I => \N__8166\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__8172\,
            I => \N__8163\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__8169\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_10\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__8166\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_10\
        );

    \I__1504\ : Odrv4
    port map (
            O => \N__8163\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_10\
        );

    \I__1503\ : InMux
    port map (
            O => \N__8156\,
            I => \N__8150\
        );

    \I__1502\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8150\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__8150\,
            I => \N__8147\
        );

    \I__1500\ : Span4Mux_v
    port map (
            O => \N__8147\,
            I => \N__8144\
        );

    \I__1499\ : Span4Mux_h
    port map (
            O => \N__8144\,
            I => \N__8141\
        );

    \I__1498\ : Sp12to4
    port map (
            O => \N__8141\,
            I => \N__8138\
        );

    \I__1497\ : Span12Mux_h
    port map (
            O => \N__8138\,
            I => \N__8135\
        );

    \I__1496\ : Odrv12
    port map (
            O => \N__8135\,
            I => miso_input_c
        );

    \I__1495\ : InMux
    port map (
            O => \N__8132\,
            I => \N__8128\
        );

    \I__1494\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8125\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__8128\,
            I => \N__8118\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__8125\,
            I => \N__8118\
        );

    \I__1491\ : InMux
    port map (
            O => \N__8124\,
            I => \N__8113\
        );

    \I__1490\ : InMux
    port map (
            O => \N__8123\,
            I => \N__8113\
        );

    \I__1489\ : Span4Mux_h
    port map (
            O => \N__8118\,
            I => \N__8110\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__8113\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_0\
        );

    \I__1487\ : Odrv4
    port map (
            O => \N__8110\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_0\
        );

    \I__1486\ : InMux
    port map (
            O => \N__8105\,
            I => \N__8102\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__8102\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_10\
        );

    \I__1484\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8096\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__8096\,
            I => \N__8093\
        );

    \I__1482\ : Span4Mux_h
    port map (
            O => \N__8093\,
            I => \N__8090\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__8090\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_15\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__8087\,
            I => \clk_out_RNI3LEM_cascade_\
        );

    \I__1479\ : CascadeMux
    port map (
            O => \N__8084\,
            I => \FSM_TEST_inst_RAPIDA.N_100_li_cascade_\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__8081\,
            I => \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5DZ0Z1_cascade_\
        );

    \I__1477\ : CEMux
    port map (
            O => \N__8078\,
            I => \N__8075\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__8075\,
            I => \N__8072\
        );

    \I__1475\ : Odrv4
    port map (
            O => \N__8072\,
            I => \N_378_i\
        );

    \I__1474\ : InMux
    port map (
            O => \N__8069\,
            I => \N__8063\
        );

    \I__1473\ : InMux
    port map (
            O => \N__8068\,
            I => \N__8063\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__8063\,
            I => \N__8058\
        );

    \I__1471\ : InMux
    port map (
            O => \N__8062\,
            I => \N__8053\
        );

    \I__1470\ : InMux
    port map (
            O => \N__8061\,
            I => \N__8053\
        );

    \I__1469\ : Span4Mux_h
    port map (
            O => \N__8058\,
            I => \N__8050\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__8053\,
            I => flag_signal
        );

    \I__1467\ : Odrv4
    port map (
            O => \N__8050\,
            I => flag_signal
        );

    \I__1466\ : InMux
    port map (
            O => \N__8045\,
            I => \N__8042\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__8042\,
            I => mosi_fast
        );

    \I__1464\ : InMux
    port map (
            O => \N__8039\,
            I => \N__8036\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__8036\,
            I => \N__8033\
        );

    \I__1462\ : Span4Mux_h
    port map (
            O => \N__8033\,
            I => \N__8030\
        );

    \I__1461\ : Odrv4
    port map (
            O => \N__8030\,
            I => mosi_slow
        );

    \I__1460\ : IoInMux
    port map (
            O => \N__8027\,
            I => \N__8024\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__8024\,
            I => \N__8021\
        );

    \I__1458\ : IoSpan4Mux
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__1457\ : Sp12to4
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__1456\ : Span12Mux_s7_h
    port map (
            O => \N__8015\,
            I => \N__8012\
        );

    \I__1455\ : Span12Mux_h
    port map (
            O => \N__8012\,
            I => \N__8009\
        );

    \I__1454\ : Span12Mux_v
    port map (
            O => \N__8009\,
            I => \N__8006\
        );

    \I__1453\ : Odrv12
    port map (
            O => \N__8006\,
            I => mosi_output_c
        );

    \I__1452\ : InMux
    port map (
            O => \N__8003\,
            I => \N__7999\
        );

    \I__1451\ : CascadeMux
    port map (
            O => \N__8002\,
            I => \N__7996\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7999\,
            I => \N__7993\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7996\,
            I => \N__7990\
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__7993\,
            I => \config_register_latched_dec_inst.DYNCNF_1Z0Z_10\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7990\,
            I => \config_register_latched_dec_inst.DYNCNF_1Z0Z_10\
        );

    \I__1446\ : IoInMux
    port map (
            O => \N__7985\,
            I => \N__7982\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7982\,
            I => \N__7979\
        );

    \I__1444\ : IoSpan4Mux
    port map (
            O => \N__7979\,
            I => \N__7976\
        );

    \I__1443\ : Sp12to4
    port map (
            O => \N__7976\,
            I => \N__7973\
        );

    \I__1442\ : Span12Mux_h
    port map (
            O => \N__7973\,
            I => \N__7970\
        );

    \I__1441\ : Odrv12
    port map (
            O => \N__7970\,
            I => s14_c
        );

    \I__1440\ : CEMux
    port map (
            O => \N__7967\,
            I => \N__7964\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__7964\,
            I => \N__7961\
        );

    \I__1438\ : Odrv12
    port map (
            O => \N__7961\,
            I => \config_register_latched_dec_inst.N_378_i_i\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7958\,
            I => \N__7955\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7955\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_64\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7952\,
            I => \N__7949\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__7949\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_65\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7946\,
            I => \N__7943\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7943\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_62\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__7940\,
            I => \N__7935\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__7939\,
            I => \N__7932\
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__7938\,
            I => \N__7910\
        );

    \I__1428\ : InMux
    port map (
            O => \N__7935\,
            I => \N__7892\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7932\,
            I => \N__7892\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7931\,
            I => \N__7892\
        );

    \I__1425\ : InMux
    port map (
            O => \N__7930\,
            I => \N__7889\
        );

    \I__1424\ : InMux
    port map (
            O => \N__7929\,
            I => \N__7882\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__7928\,
            I => \N__7872\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__7927\,
            I => \N__7869\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__7926\,
            I => \N__7866\
        );

    \I__1420\ : CascadeMux
    port map (
            O => \N__7925\,
            I => \N__7860\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__7924\,
            I => \N__7855\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__7923\,
            I => \N__7852\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__7922\,
            I => \N__7845\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__7921\,
            I => \N__7842\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__7920\,
            I => \N__7838\
        );

    \I__1414\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7824\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__7918\,
            I => \N__7821\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__7917\,
            I => \N__7818\
        );

    \I__1411\ : CascadeMux
    port map (
            O => \N__7916\,
            I => \N__7815\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__7915\,
            I => \N__7808\
        );

    \I__1409\ : CascadeMux
    port map (
            O => \N__7914\,
            I => \N__7804\
        );

    \I__1408\ : CascadeMux
    port map (
            O => \N__7913\,
            I => \N__7801\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7791\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7791\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7786\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7907\,
            I => \N__7786\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__7906\,
            I => \N__7782\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__7905\,
            I => \N__7778\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__7904\,
            I => \N__7775\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__7903\,
            I => \N__7770\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__7902\,
            I => \N__7767\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__7901\,
            I => \N__7763\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__7900\,
            I => \N__7758\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__7899\,
            I => \N__7754\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__7892\,
            I => \N__7749\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__7889\,
            I => \N__7746\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7888\,
            I => \N__7743\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7887\,
            I => \N__7736\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7886\,
            I => \N__7736\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7885\,
            I => \N__7736\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__7882\,
            I => \N__7733\
        );

    \I__1388\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7722\
        );

    \I__1387\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7722\
        );

    \I__1386\ : InMux
    port map (
            O => \N__7879\,
            I => \N__7722\
        );

    \I__1385\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7722\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7722\
        );

    \I__1383\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7707\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7707\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7872\,
            I => \N__7707\
        );

    \I__1380\ : InMux
    port map (
            O => \N__7869\,
            I => \N__7707\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7866\,
            I => \N__7707\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7865\,
            I => \N__7707\
        );

    \I__1377\ : InMux
    port map (
            O => \N__7864\,
            I => \N__7707\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7863\,
            I => \N__7700\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7860\,
            I => \N__7700\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7859\,
            I => \N__7700\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7858\,
            I => \N__7691\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7855\,
            I => \N__7691\
        );

    \I__1371\ : InMux
    port map (
            O => \N__7852\,
            I => \N__7691\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7851\,
            I => \N__7691\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7850\,
            I => \N__7688\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7849\,
            I => \N__7685\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7848\,
            I => \N__7682\
        );

    \I__1366\ : InMux
    port map (
            O => \N__7845\,
            I => \N__7671\
        );

    \I__1365\ : InMux
    port map (
            O => \N__7842\,
            I => \N__7671\
        );

    \I__1364\ : InMux
    port map (
            O => \N__7841\,
            I => \N__7671\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7838\,
            I => \N__7671\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7837\,
            I => \N__7671\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7836\,
            I => \N__7654\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7835\,
            I => \N__7654\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7834\,
            I => \N__7654\
        );

    \I__1358\ : InMux
    port map (
            O => \N__7833\,
            I => \N__7654\
        );

    \I__1357\ : InMux
    port map (
            O => \N__7832\,
            I => \N__7645\
        );

    \I__1356\ : InMux
    port map (
            O => \N__7831\,
            I => \N__7645\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7830\,
            I => \N__7645\
        );

    \I__1354\ : InMux
    port map (
            O => \N__7829\,
            I => \N__7645\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__7828\,
            I => \N__7641\
        );

    \I__1352\ : InMux
    port map (
            O => \N__7827\,
            I => \N__7635\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7824\,
            I => \N__7632\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7821\,
            I => \N__7621\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7818\,
            I => \N__7621\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7815\,
            I => \N__7621\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7814\,
            I => \N__7621\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7813\,
            I => \N__7621\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7617\
        );

    \I__1344\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7614\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7808\,
            I => \N__7609\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7807\,
            I => \N__7609\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7804\,
            I => \N__7602\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7801\,
            I => \N__7602\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7800\,
            I => \N__7602\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7799\,
            I => \N__7593\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7798\,
            I => \N__7593\
        );

    \I__1336\ : InMux
    port map (
            O => \N__7797\,
            I => \N__7593\
        );

    \I__1335\ : InMux
    port map (
            O => \N__7796\,
            I => \N__7593\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7791\,
            I => \N__7588\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__7786\,
            I => \N__7588\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7785\,
            I => \N__7573\
        );

    \I__1331\ : InMux
    port map (
            O => \N__7782\,
            I => \N__7573\
        );

    \I__1330\ : InMux
    port map (
            O => \N__7781\,
            I => \N__7573\
        );

    \I__1329\ : InMux
    port map (
            O => \N__7778\,
            I => \N__7573\
        );

    \I__1328\ : InMux
    port map (
            O => \N__7775\,
            I => \N__7573\
        );

    \I__1327\ : InMux
    port map (
            O => \N__7774\,
            I => \N__7573\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7773\,
            I => \N__7573\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7770\,
            I => \N__7548\
        );

    \I__1324\ : InMux
    port map (
            O => \N__7767\,
            I => \N__7548\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7766\,
            I => \N__7548\
        );

    \I__1322\ : InMux
    port map (
            O => \N__7763\,
            I => \N__7548\
        );

    \I__1321\ : InMux
    port map (
            O => \N__7762\,
            I => \N__7548\
        );

    \I__1320\ : InMux
    port map (
            O => \N__7761\,
            I => \N__7548\
        );

    \I__1319\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7537\
        );

    \I__1318\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7537\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7754\,
            I => \N__7537\
        );

    \I__1316\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7537\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7752\,
            I => \N__7537\
        );

    \I__1314\ : Span4Mux_v
    port map (
            O => \N__7749\,
            I => \N__7525\
        );

    \I__1313\ : Span4Mux_v
    port map (
            O => \N__7746\,
            I => \N__7525\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__7743\,
            I => \N__7525\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__7736\,
            I => \N__7525\
        );

    \I__1310\ : Span4Mux_v
    port map (
            O => \N__7733\,
            I => \N__7514\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__7722\,
            I => \N__7514\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__7707\,
            I => \N__7514\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__7700\,
            I => \N__7514\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__7691\,
            I => \N__7514\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__7688\,
            I => \N__7509\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__7685\,
            I => \N__7509\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__7682\,
            I => \N__7504\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__7671\,
            I => \N__7504\
        );

    \I__1301\ : InMux
    port map (
            O => \N__7670\,
            I => \N__7487\
        );

    \I__1300\ : InMux
    port map (
            O => \N__7669\,
            I => \N__7487\
        );

    \I__1299\ : InMux
    port map (
            O => \N__7668\,
            I => \N__7487\
        );

    \I__1298\ : InMux
    port map (
            O => \N__7667\,
            I => \N__7487\
        );

    \I__1297\ : InMux
    port map (
            O => \N__7666\,
            I => \N__7487\
        );

    \I__1296\ : InMux
    port map (
            O => \N__7665\,
            I => \N__7487\
        );

    \I__1295\ : InMux
    port map (
            O => \N__7664\,
            I => \N__7487\
        );

    \I__1294\ : InMux
    port map (
            O => \N__7663\,
            I => \N__7487\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__7654\,
            I => \N__7482\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__7645\,
            I => \N__7482\
        );

    \I__1291\ : InMux
    port map (
            O => \N__7644\,
            I => \N__7471\
        );

    \I__1290\ : InMux
    port map (
            O => \N__7641\,
            I => \N__7471\
        );

    \I__1289\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7471\
        );

    \I__1288\ : InMux
    port map (
            O => \N__7639\,
            I => \N__7471\
        );

    \I__1287\ : InMux
    port map (
            O => \N__7638\,
            I => \N__7471\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__7635\,
            I => \N__7468\
        );

    \I__1285\ : Span4Mux_h
    port map (
            O => \N__7632\,
            I => \N__7463\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__7621\,
            I => \N__7463\
        );

    \I__1283\ : InMux
    port map (
            O => \N__7620\,
            I => \N__7460\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__7617\,
            I => \N__7454\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__7614\,
            I => \N__7447\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__7609\,
            I => \N__7447\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__7602\,
            I => \N__7447\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__7593\,
            I => \N__7444\
        );

    \I__1277\ : Span4Mux_h
    port map (
            O => \N__7588\,
            I => \N__7439\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__7573\,
            I => \N__7439\
        );

    \I__1275\ : InMux
    port map (
            O => \N__7572\,
            I => \N__7432\
        );

    \I__1274\ : InMux
    port map (
            O => \N__7571\,
            I => \N__7432\
        );

    \I__1273\ : InMux
    port map (
            O => \N__7570\,
            I => \N__7432\
        );

    \I__1272\ : InMux
    port map (
            O => \N__7569\,
            I => \N__7427\
        );

    \I__1271\ : InMux
    port map (
            O => \N__7568\,
            I => \N__7427\
        );

    \I__1270\ : InMux
    port map (
            O => \N__7567\,
            I => \N__7420\
        );

    \I__1269\ : InMux
    port map (
            O => \N__7566\,
            I => \N__7420\
        );

    \I__1268\ : InMux
    port map (
            O => \N__7565\,
            I => \N__7420\
        );

    \I__1267\ : InMux
    port map (
            O => \N__7564\,
            I => \N__7411\
        );

    \I__1266\ : InMux
    port map (
            O => \N__7563\,
            I => \N__7411\
        );

    \I__1265\ : InMux
    port map (
            O => \N__7562\,
            I => \N__7411\
        );

    \I__1264\ : InMux
    port map (
            O => \N__7561\,
            I => \N__7411\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__7548\,
            I => \N__7406\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__7537\,
            I => \N__7406\
        );

    \I__1261\ : InMux
    port map (
            O => \N__7536\,
            I => \N__7399\
        );

    \I__1260\ : InMux
    port map (
            O => \N__7535\,
            I => \N__7399\
        );

    \I__1259\ : InMux
    port map (
            O => \N__7534\,
            I => \N__7399\
        );

    \I__1258\ : Span4Mux_h
    port map (
            O => \N__7525\,
            I => \N__7392\
        );

    \I__1257\ : Span4Mux_v
    port map (
            O => \N__7514\,
            I => \N__7392\
        );

    \I__1256\ : Span4Mux_v
    port map (
            O => \N__7509\,
            I => \N__7392\
        );

    \I__1255\ : Span4Mux_v
    port map (
            O => \N__7504\,
            I => \N__7383\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__7487\,
            I => \N__7383\
        );

    \I__1253\ : Span4Mux_v
    port map (
            O => \N__7482\,
            I => \N__7383\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__7471\,
            I => \N__7383\
        );

    \I__1251\ : Span4Mux_v
    port map (
            O => \N__7468\,
            I => \N__7376\
        );

    \I__1250\ : Span4Mux_h
    port map (
            O => \N__7463\,
            I => \N__7376\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__7460\,
            I => \N__7376\
        );

    \I__1248\ : InMux
    port map (
            O => \N__7459\,
            I => \N__7369\
        );

    \I__1247\ : InMux
    port map (
            O => \N__7458\,
            I => \N__7369\
        );

    \I__1246\ : InMux
    port map (
            O => \N__7457\,
            I => \N__7369\
        );

    \I__1245\ : Odrv12
    port map (
            O => \N__7454\,
            I => \FSM_TEST_inst_slow.current_stateZ0Z_1\
        );

    \I__1244\ : Odrv12
    port map (
            O => \N__7447\,
            I => \FSM_TEST_inst_slow.current_stateZ0Z_1\
        );

    \I__1243\ : Odrv4
    port map (
            O => \N__7444\,
            I => \FSM_TEST_inst_slow.current_stateZ0Z_1\
        );

    \I__1242\ : Odrv4
    port map (
            O => \N__7439\,
            I => \FSM_TEST_inst_slow.current_stateZ0Z_1\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__7432\,
            I => \FSM_TEST_inst_slow.current_stateZ0Z_1\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__7427\,
            I => \FSM_TEST_inst_slow.current_stateZ0Z_1\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__7420\,
            I => \FSM_TEST_inst_slow.current_stateZ0Z_1\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__7411\,
            I => \FSM_TEST_inst_slow.current_stateZ0Z_1\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__7406\,
            I => \FSM_TEST_inst_slow.current_stateZ0Z_1\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__7399\,
            I => \FSM_TEST_inst_slow.current_stateZ0Z_1\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__7392\,
            I => \FSM_TEST_inst_slow.current_stateZ0Z_1\
        );

    \I__1234\ : Odrv4
    port map (
            O => \N__7383\,
            I => \FSM_TEST_inst_slow.current_stateZ0Z_1\
        );

    \I__1233\ : Odrv4
    port map (
            O => \N__7376\,
            I => \FSM_TEST_inst_slow.current_stateZ0Z_1\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__7369\,
            I => \FSM_TEST_inst_slow.current_stateZ0Z_1\
        );

    \I__1231\ : InMux
    port map (
            O => \N__7340\,
            I => \N__7337\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__7337\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_63\
        );

    \I__1229\ : CEMux
    port map (
            O => \N__7334\,
            I => \N__7259\
        );

    \I__1228\ : CEMux
    port map (
            O => \N__7333\,
            I => \N__7259\
        );

    \I__1227\ : CEMux
    port map (
            O => \N__7332\,
            I => \N__7259\
        );

    \I__1226\ : CEMux
    port map (
            O => \N__7331\,
            I => \N__7259\
        );

    \I__1225\ : CEMux
    port map (
            O => \N__7330\,
            I => \N__7259\
        );

    \I__1224\ : CEMux
    port map (
            O => \N__7329\,
            I => \N__7259\
        );

    \I__1223\ : CEMux
    port map (
            O => \N__7328\,
            I => \N__7259\
        );

    \I__1222\ : CEMux
    port map (
            O => \N__7327\,
            I => \N__7259\
        );

    \I__1221\ : CEMux
    port map (
            O => \N__7326\,
            I => \N__7259\
        );

    \I__1220\ : CEMux
    port map (
            O => \N__7325\,
            I => \N__7259\
        );

    \I__1219\ : CEMux
    port map (
            O => \N__7324\,
            I => \N__7259\
        );

    \I__1218\ : CEMux
    port map (
            O => \N__7323\,
            I => \N__7259\
        );

    \I__1217\ : CEMux
    port map (
            O => \N__7322\,
            I => \N__7259\
        );

    \I__1216\ : CEMux
    port map (
            O => \N__7321\,
            I => \N__7259\
        );

    \I__1215\ : CEMux
    port map (
            O => \N__7320\,
            I => \N__7259\
        );

    \I__1214\ : CEMux
    port map (
            O => \N__7319\,
            I => \N__7259\
        );

    \I__1213\ : CEMux
    port map (
            O => \N__7318\,
            I => \N__7259\
        );

    \I__1212\ : CEMux
    port map (
            O => \N__7317\,
            I => \N__7259\
        );

    \I__1211\ : CEMux
    port map (
            O => \N__7316\,
            I => \N__7259\
        );

    \I__1210\ : CEMux
    port map (
            O => \N__7315\,
            I => \N__7259\
        );

    \I__1209\ : CEMux
    port map (
            O => \N__7314\,
            I => \N__7259\
        );

    \I__1208\ : CEMux
    port map (
            O => \N__7313\,
            I => \N__7259\
        );

    \I__1207\ : CEMux
    port map (
            O => \N__7312\,
            I => \N__7259\
        );

    \I__1206\ : CEMux
    port map (
            O => \N__7311\,
            I => \N__7259\
        );

    \I__1205\ : CEMux
    port map (
            O => \N__7310\,
            I => \N__7259\
        );

    \I__1204\ : GlobalMux
    port map (
            O => \N__7259\,
            I => \N__7256\
        );

    \I__1203\ : gio2CtrlBuf
    port map (
            O => \N__7256\,
            I => \FSM_TEST_inst_slow.N_374_g\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__7253\,
            I => \counter_RNIFD27_2_cascade_\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__7250\,
            I => \N_3_0_cascade_\
        );

    \I__1200\ : InMux
    port map (
            O => \N__7247\,
            I => \N__7244\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__7244\,
            I => \N_2_0\
        );

    \I__1198\ : CEMux
    port map (
            O => \N__7241\,
            I => \N__7235\
        );

    \I__1197\ : InMux
    port map (
            O => \N__7240\,
            I => \N__7228\
        );

    \I__1196\ : InMux
    port map (
            O => \N__7239\,
            I => \N__7228\
        );

    \I__1195\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7228\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__7235\,
            I => \N__7222\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__7228\,
            I => \N__7219\
        );

    \I__1192\ : InMux
    port map (
            O => \N__7227\,
            I => \N__7212\
        );

    \I__1191\ : InMux
    port map (
            O => \N__7226\,
            I => \N__7212\
        );

    \I__1190\ : InMux
    port map (
            O => \N__7225\,
            I => \N__7212\
        );

    \I__1189\ : Span4Mux_h
    port map (
            O => \N__7222\,
            I => \N__7205\
        );

    \I__1188\ : Span4Mux_v
    port map (
            O => \N__7219\,
            I => \N__7200\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__7212\,
            I => \N__7200\
        );

    \I__1186\ : InMux
    port map (
            O => \N__7211\,
            I => \N__7191\
        );

    \I__1185\ : InMux
    port map (
            O => \N__7210\,
            I => \N__7191\
        );

    \I__1184\ : InMux
    port map (
            O => \N__7209\,
            I => \N__7191\
        );

    \I__1183\ : InMux
    port map (
            O => \N__7208\,
            I => \N__7191\
        );

    \I__1182\ : Odrv4
    port map (
            O => \N__7205\,
            I => \counter_RNISR1F_2\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__7200\,
            I => \counter_RNISR1F_2\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__7191\,
            I => \counter_RNISR1F_2\
        );

    \I__1179\ : InMux
    port map (
            O => \N__7184\,
            I => \N__7181\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__7181\,
            I => \FSM_TEST_inst_RAPIDA.CLK_uC_3Z0Z_0\
        );

    \I__1177\ : InMux
    port map (
            O => \N__7178\,
            I => \N__7175\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__7175\,
            I => \FSM_TEST_inst_RAPIDA.CLK_uC_4Z0Z_0\
        );

    \I__1175\ : InMux
    port map (
            O => \N__7172\,
            I => \N__7169\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__7169\,
            I => \FSM_TEST_inst_RAPIDA.CLK_uC_5Z0Z_0\
        );

    \I__1173\ : InMux
    port map (
            O => \N__7166\,
            I => \N__7163\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__7163\,
            I => \FSM_TEST_inst_RAPIDA.CLK_uC_6Z0Z_0\
        );

    \I__1171\ : InMux
    port map (
            O => \N__7160\,
            I => \N__7157\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__7157\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_57\
        );

    \I__1169\ : InMux
    port map (
            O => \N__7154\,
            I => \N__7151\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__7151\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_60\
        );

    \I__1167\ : InMux
    port map (
            O => \N__7148\,
            I => \N__7145\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__7145\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_58\
        );

    \I__1165\ : InMux
    port map (
            O => \N__7142\,
            I => \N__7139\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__7139\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_59\
        );

    \I__1163\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7133\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__7133\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_61\
        );

    \I__1161\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7127\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__7127\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_66\
        );

    \I__1159\ : InMux
    port map (
            O => \N__7124\,
            I => \N__7121\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__7121\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_13\
        );

    \I__1157\ : InMux
    port map (
            O => \N__7118\,
            I => \N__7115\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__7115\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_14\
        );

    \I__1155\ : InMux
    port map (
            O => \N__7112\,
            I => \N__7109\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__7109\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_18\
        );

    \I__1153\ : InMux
    port map (
            O => \N__7106\,
            I => \N__7103\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__7103\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_24\
        );

    \I__1151\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7097\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__7097\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_78\
        );

    \I__1149\ : InMux
    port map (
            O => \N__7094\,
            I => \N__7091\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__7091\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_77\
        );

    \I__1147\ : InMux
    port map (
            O => \N__7088\,
            I => \N__7085\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__7085\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_25\
        );

    \I__1145\ : InMux
    port map (
            O => \N__7082\,
            I => \N__7079\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__7079\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_26\
        );

    \I__1143\ : InMux
    port map (
            O => \N__7076\,
            I => \N__7073\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__7073\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_0\
        );

    \I__1141\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7067\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__7067\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_1\
        );

    \I__1139\ : InMux
    port map (
            O => \N__7064\,
            I => \N__7061\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__7061\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_4\
        );

    \I__1137\ : InMux
    port map (
            O => \N__7058\,
            I => \N__7055\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__7055\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_5\
        );

    \I__1135\ : InMux
    port map (
            O => \N__7052\,
            I => \N__7049\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__7049\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_2\
        );

    \I__1133\ : InMux
    port map (
            O => \N__7046\,
            I => \N__7043\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__7043\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_3\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__7040\,
            I => \FSM_TEST_inst_RAPIDA.counter_din_3_i_0_2_cascade_\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__7037\,
            I => \FSM_TEST_inst_RAPIDA.G_24_0_o4_2_cascade_\
        );

    \I__1129\ : InMux
    port map (
            O => \N__7034\,
            I => \N__7031\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__7031\,
            I => \N__7028\
        );

    \I__1127\ : Odrv4
    port map (
            O => \N__7028\,
            I => \FSM_TEST_inst_RAPIDA.G_24_0_a4_0_1\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__7025\,
            I => \N__7022\
        );

    \I__1125\ : InMux
    port map (
            O => \N__7022\,
            I => \N__7018\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__7021\,
            I => \N__7014\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__7018\,
            I => \N__7011\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__7017\,
            I => \N__7008\
        );

    \I__1121\ : InMux
    port map (
            O => \N__7014\,
            I => \N__7005\
        );

    \I__1120\ : Span4Mux_h
    port map (
            O => \N__7011\,
            I => \N__7002\
        );

    \I__1119\ : InMux
    port map (
            O => \N__7008\,
            I => \N__6999\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__7005\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_6\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__7002\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_6\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6999\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_6\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6992\,
            I => \N__6989\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6989\,
            I => \N__6986\
        );

    \I__1113\ : Span4Mux_h
    port map (
            O => \N__6986\,
            I => \N__6980\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6985\,
            I => \N__6977\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6984\,
            I => \N__6972\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6983\,
            I => \N__6972\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__6980\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_3\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6977\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_3\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6972\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_3\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6965\,
            I => \N__6962\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__6962\,
            I => \FSM_TEST_inst_RAPIDA.G_24_0_a4_0_5\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6959\,
            I => \N__6956\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__6956\,
            I => \FSM_TEST_inst_RAPIDA.N_18_0\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__6953\,
            I => \FSM_TEST_inst_RAPIDA.G_24_0_a4_0_6_cascade_\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6950\,
            I => \N__6947\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6947\,
            I => \FSM_TEST_inst_RAPIDA.N_9_1\
        );

    \I__1099\ : InMux
    port map (
            O => \N__6944\,
            I => \N__6937\
        );

    \I__1098\ : InMux
    port map (
            O => \N__6943\,
            I => \N__6937\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__6942\,
            I => \N__6934\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__6937\,
            I => \N__6931\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6934\,
            I => \N__6928\
        );

    \I__1094\ : Span4Mux_v
    port map (
            O => \N__6931\,
            I => \N__6925\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6928\,
            I => \FSM_TEST_inst_slow.counter_dinZ0Z_3\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__6925\,
            I => \FSM_TEST_inst_slow.counter_dinZ0Z_3\
        );

    \I__1091\ : InMux
    port map (
            O => \N__6920\,
            I => \N__6917\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__6917\,
            I => \N__6913\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__6916\,
            I => \N__6909\
        );

    \I__1088\ : Span4Mux_h
    port map (
            O => \N__6913\,
            I => \N__6905\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6912\,
            I => \N__6898\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6909\,
            I => \N__6898\
        );

    \I__1085\ : InMux
    port map (
            O => \N__6908\,
            I => \N__6898\
        );

    \I__1084\ : Odrv4
    port map (
            O => \N__6905\,
            I => \FSM_TEST_inst_slow.counter_dinZ0Z_2\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__6898\,
            I => \FSM_TEST_inst_slow.counter_dinZ0Z_2\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6884\
        );

    \I__1081\ : InMux
    port map (
            O => \N__6892\,
            I => \N__6884\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6891\,
            I => \N__6884\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6884\,
            I => \N__6881\
        );

    \I__1078\ : Span4Mux_v
    port map (
            O => \N__6881\,
            I => \N__6878\
        );

    \I__1077\ : Odrv4
    port map (
            O => \N__6878\,
            I => \FSM_TEST_inst_slow.N_106_0\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__6875\,
            I => \FSM_TEST_inst_slow.current_state_RNO_8Z0Z_0_cascade_\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6872\,
            I => \N__6869\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__6869\,
            I => \FSM_TEST_inst_slow.current_state_RNO_1Z0Z_0\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6866\,
            I => \N__6863\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__6863\,
            I => \N__6860\
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__6860\,
            I => \FSM_TEST_inst_slow.N_134\
        );

    \I__1070\ : CascadeMux
    port map (
            O => \N__6857\,
            I => \FSM_TEST_inst_slow.current_state_RNO_2Z0Z_0_cascade_\
        );

    \I__1069\ : IoInMux
    port map (
            O => \N__6854\,
            I => \N__6851\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6851\,
            I => \N__6848\
        );

    \I__1067\ : Span4Mux_s1_v
    port map (
            O => \N__6848\,
            I => \N__6845\
        );

    \I__1066\ : Sp12to4
    port map (
            O => \N__6845\,
            I => \N__6842\
        );

    \I__1065\ : Span12Mux_s11_h
    port map (
            O => \N__6842\,
            I => \N__6839\
        );

    \I__1064\ : Span12Mux_v
    port map (
            O => \N__6839\,
            I => \N__6836\
        );

    \I__1063\ : Odrv12
    port map (
            O => \N__6836\,
            I => s12_c
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__6833\,
            I => \N__6829\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6832\,
            I => \N__6824\
        );

    \I__1060\ : InMux
    port map (
            O => \N__6829\,
            I => \N__6824\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6824\,
            I => \config_register_latched_dec_inst.DYNCNF_1Z0Z_8\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6821\,
            I => \N__6815\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6820\,
            I => \N__6815\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6815\,
            I => \config_register_latched_dec_inst.DYNCNF_1Z0Z_9\
        );

    \I__1055\ : IoInMux
    port map (
            O => \N__6812\,
            I => \N__6809\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__6809\,
            I => \N__6806\
        );

    \I__1053\ : Span12Mux_s11_h
    port map (
            O => \N__6806\,
            I => \N__6803\
        );

    \I__1052\ : Odrv12
    port map (
            O => \N__6803\,
            I => s13_c
        );

    \I__1051\ : InMux
    port map (
            O => \N__6800\,
            I => \N__6794\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6799\,
            I => \N__6794\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6794\,
            I => \config_register_latched_dec_inst.DYNCNF_1Z0Z_0\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6788\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__6788\,
            I => \N__6785\
        );

    \I__1046\ : Span4Mux_h
    port map (
            O => \N__6785\,
            I => \N__6782\
        );

    \I__1045\ : Span4Mux_v
    port map (
            O => \N__6782\,
            I => \N__6779\
        );

    \I__1044\ : Sp12to4
    port map (
            O => \N__6779\,
            I => \N__6776\
        );

    \I__1043\ : Span12Mux_v
    port map (
            O => \N__6776\,
            I => \N__6773\
        );

    \I__1042\ : Odrv12
    port map (
            O => \N__6773\,
            I => \config_register_latched_dec_inst.DYNCNF_0\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6770\,
            I => \N__6767\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6767\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_6\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6764\,
            I => \N__6761\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__6761\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_56\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6758\,
            I => \N__6755\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6755\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_69\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6752\,
            I => \N__6749\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6749\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_68\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6746\,
            I => \N__6743\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6743\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_67\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__6740\,
            I => \FSM_TEST_inst_slow.N_108_li_cascade_\
        );

    \I__1030\ : IoInMux
    port map (
            O => \N__6737\,
            I => \N__6734\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6734\,
            I => \N__6731\
        );

    \I__1028\ : Span12Mux_s5_h
    port map (
            O => \N__6731\,
            I => \N__6728\
        );

    \I__1027\ : Odrv12
    port map (
            O => \N__6728\,
            I => \FSM_TEST_inst_slow.current_state_RNIR2L81_0Z0Z_1\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6725\,
            I => \N__6722\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__6722\,
            I => \FSM_TEST_inst_slow.current_state_cnv_0_1\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6719\,
            I => \N__6709\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6718\,
            I => \N__6709\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6717\,
            I => \N__6709\
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__6716\,
            I => \N__6706\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__6709\,
            I => \N__6703\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6706\,
            I => \N__6700\
        );

    \I__1018\ : Span4Mux_h
    port map (
            O => \N__6703\,
            I => \N__6697\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__6700\,
            I => \FSM_TEST_inst_slow.N_108_li\
        );

    \I__1016\ : Odrv4
    port map (
            O => \N__6697\,
            I => \FSM_TEST_inst_slow.N_108_li\
        );

    \I__1015\ : InMux
    port map (
            O => \N__6692\,
            I => \N__6689\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__6689\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_7\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6686\,
            I => \N__6683\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6683\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_8\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6677\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__6677\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_9\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6671\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6671\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_53\
        );

    \I__1007\ : InMux
    port map (
            O => \N__6668\,
            I => \N__6665\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6665\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_10\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6662\,
            I => \N__6659\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__6659\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_11\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6656\,
            I => \N__6653\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6653\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_54\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6650\,
            I => \N__6647\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__6647\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_55\
        );

    \I__999\ : InMux
    port map (
            O => \N__6644\,
            I => \N__6641\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__6641\,
            I => \N__6638\
        );

    \I__997\ : Odrv12
    port map (
            O => \N__6638\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_50\
        );

    \I__996\ : InMux
    port map (
            O => \N__6635\,
            I => \N__6632\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__6632\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_51\
        );

    \I__994\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6626\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__6626\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_5\
        );

    \I__992\ : InMux
    port map (
            O => \N__6623\,
            I => \N__6620\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__6620\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_23\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__6617\,
            I => \N__6613\
        );

    \I__989\ : InMux
    port map (
            O => \N__6616\,
            I => \N__6610\
        );

    \I__988\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6606\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__6610\,
            I => \N__6603\
        );

    \I__986\ : InMux
    port map (
            O => \N__6609\,
            I => \N__6599\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__6606\,
            I => \N__6596\
        );

    \I__984\ : Span4Mux_v
    port map (
            O => \N__6603\,
            I => \N__6593\
        );

    \I__983\ : InMux
    port map (
            O => \N__6602\,
            I => \N__6590\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__6599\,
            I => \N__6587\
        );

    \I__981\ : Odrv12
    port map (
            O => \N__6596\,
            I => \CONSTANT_ONE_NET\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__6593\,
            I => \CONSTANT_ONE_NET\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__6590\,
            I => \CONSTANT_ONE_NET\
        );

    \I__978\ : Odrv4
    port map (
            O => \N__6587\,
            I => \CONSTANT_ONE_NET\
        );

    \I__977\ : InMux
    port map (
            O => \N__6578\,
            I => \N__6575\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__6575\,
            I => \N__6572\
        );

    \I__975\ : Odrv4
    port map (
            O => \N__6572\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_86\
        );

    \I__974\ : InMux
    port map (
            O => \N__6569\,
            I => \N__6566\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__6566\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_84\
        );

    \I__972\ : InMux
    port map (
            O => \N__6563\,
            I => \N__6560\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__6560\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_85\
        );

    \I__970\ : InMux
    port map (
            O => \N__6557\,
            I => \N__6554\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__6554\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_82\
        );

    \I__968\ : InMux
    port map (
            O => \N__6551\,
            I => \N__6548\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__6548\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_83\
        );

    \I__966\ : InMux
    port map (
            O => \N__6545\,
            I => \N__6542\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__6542\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_12\
        );

    \I__964\ : InMux
    port map (
            O => \N__6539\,
            I => \N__6536\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__6536\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_52\
        );

    \I__962\ : CascadeMux
    port map (
            O => \N__6533\,
            I => \FSM_TEST_inst_RAPIDA.counter_idlelde_2_cascade_\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__6530\,
            I => \N__6525\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__6529\,
            I => \N__6522\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__6528\,
            I => \N__6517\
        );

    \I__958\ : InMux
    port map (
            O => \N__6525\,
            I => \N__6510\
        );

    \I__957\ : InMux
    port map (
            O => \N__6522\,
            I => \N__6510\
        );

    \I__956\ : InMux
    port map (
            O => \N__6521\,
            I => \N__6510\
        );

    \I__955\ : InMux
    port map (
            O => \N__6520\,
            I => \N__6507\
        );

    \I__954\ : InMux
    port map (
            O => \N__6517\,
            I => \N__6504\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__6510\,
            I => \N__6501\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__6507\,
            I => \N__6498\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__6504\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1\
        );

    \I__950\ : Odrv4
    port map (
            O => \N__6501\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1\
        );

    \I__949\ : Odrv4
    port map (
            O => \N__6498\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1\
        );

    \I__948\ : CascadeMux
    port map (
            O => \N__6491\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1_cascade_\
        );

    \I__947\ : InMux
    port map (
            O => \N__6488\,
            I => \N__6475\
        );

    \I__946\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6475\
        );

    \I__945\ : InMux
    port map (
            O => \N__6486\,
            I => \N__6475\
        );

    \I__944\ : InMux
    port map (
            O => \N__6485\,
            I => \N__6475\
        );

    \I__943\ : InMux
    port map (
            O => \N__6484\,
            I => \N__6472\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__6475\,
            I => \N__6467\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__6472\,
            I => \N__6467\
        );

    \I__940\ : Span4Mux_h
    port map (
            O => \N__6467\,
            I => \N__6464\
        );

    \I__939\ : Odrv4
    port map (
            O => \N__6464\,
            I => \FSM_TEST_inst_RAPIDA.N_126_1_i\
        );

    \I__938\ : InMux
    port map (
            O => \N__6461\,
            I => \N__6456\
        );

    \I__937\ : InMux
    port map (
            O => \N__6460\,
            I => \N__6453\
        );

    \I__936\ : InMux
    port map (
            O => \N__6459\,
            I => \N__6450\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__6456\,
            I => \N__6445\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__6453\,
            I => \N__6445\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__6450\,
            I => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_1\
        );

    \I__932\ : Odrv4
    port map (
            O => \N__6445\,
            I => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_1\
        );

    \I__931\ : CascadeMux
    port map (
            O => \N__6440\,
            I => \N__6435\
        );

    \I__930\ : InMux
    port map (
            O => \N__6439\,
            I => \N__6431\
        );

    \I__929\ : InMux
    port map (
            O => \N__6438\,
            I => \N__6424\
        );

    \I__928\ : InMux
    port map (
            O => \N__6435\,
            I => \N__6424\
        );

    \I__927\ : InMux
    port map (
            O => \N__6434\,
            I => \N__6424\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__6431\,
            I => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_2\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__6424\,
            I => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_2\
        );

    \I__924\ : InMux
    port map (
            O => \N__6419\,
            I => \N__6412\
        );

    \I__923\ : InMux
    port map (
            O => \N__6418\,
            I => \N__6412\
        );

    \I__922\ : InMux
    port map (
            O => \N__6417\,
            I => \N__6409\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__6412\,
            I => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_0\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__6409\,
            I => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_0\
        );

    \I__919\ : InMux
    port map (
            O => \N__6404\,
            I => \N__6401\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__6401\,
            I => \FSM_TEST_inst_RAPIDA.G_24_0_a4_1_5\
        );

    \I__917\ : InMux
    port map (
            O => \N__6398\,
            I => \N__6395\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__6395\,
            I => \N__6392\
        );

    \I__915\ : Odrv4
    port map (
            O => \N__6392\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_6\
        );

    \I__914\ : InMux
    port map (
            O => \N__6389\,
            I => \N__6386\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__6386\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_19\
        );

    \I__912\ : InMux
    port map (
            O => \N__6383\,
            I => \N__6380\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__6380\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_20\
        );

    \I__910\ : InMux
    port map (
            O => \N__6377\,
            I => \N__6374\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__6374\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_21\
        );

    \I__908\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6368\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__6368\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_22\
        );

    \I__906\ : InMux
    port map (
            O => \N__6365\,
            I => \N__6362\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__6362\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_3\
        );

    \I__904\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6356\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__6356\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_4\
        );

    \I__902\ : InMux
    port map (
            O => \N__6353\,
            I => \N__6350\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__6350\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_5\
        );

    \I__900\ : InMux
    port map (
            O => \N__6347\,
            I => \N__6344\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__6344\,
            I => \FSM_TEST_inst_RAPIDA.counter_idle_cry_3_THRU_CO\
        );

    \I__898\ : InMux
    port map (
            O => \N__6341\,
            I => \N__6338\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__6338\,
            I => \FSM_TEST_inst_RAPIDA.flag_input_regZ0\
        );

    \I__896\ : InMux
    port map (
            O => \N__6335\,
            I => \N__6332\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__6332\,
            I => \FSM_TEST_inst_RAPIDA.G_24_0_a4_1_4\
        );

    \I__894\ : InMux
    port map (
            O => \N__6329\,
            I => \N__6326\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__6326\,
            I => \FSM_TEST_inst_RAPIDA.counter_idle_cry_1_THRU_CO\
        );

    \I__892\ : InMux
    port map (
            O => \N__6323\,
            I => \N__6320\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__6320\,
            I => \FSM_TEST_inst_RAPIDA.counter_idle_cry_2_THRU_CO\
        );

    \I__890\ : InMux
    port map (
            O => \N__6317\,
            I => \N__6311\
        );

    \I__889\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6304\
        );

    \I__888\ : InMux
    port map (
            O => \N__6315\,
            I => \N__6304\
        );

    \I__887\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6304\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__6311\,
            I => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_4\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__6304\,
            I => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_4\
        );

    \I__884\ : CascadeMux
    port map (
            O => \N__6299\,
            I => \N__6295\
        );

    \I__883\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6290\
        );

    \I__882\ : InMux
    port map (
            O => \N__6295\,
            I => \N__6283\
        );

    \I__881\ : InMux
    port map (
            O => \N__6294\,
            I => \N__6283\
        );

    \I__880\ : InMux
    port map (
            O => \N__6293\,
            I => \N__6283\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__6290\,
            I => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_3\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__6283\,
            I => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_3\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__6278\,
            I => \N__6273\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__6277\,
            I => \N__6270\
        );

    \I__875\ : InMux
    port map (
            O => \N__6276\,
            I => \N__6267\
        );

    \I__874\ : InMux
    port map (
            O => \N__6273\,
            I => \N__6264\
        );

    \I__873\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6261\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__6267\,
            I => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_5\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__6264\,
            I => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_5\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__6261\,
            I => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_5\
        );

    \I__869\ : InMux
    port map (
            O => \N__6254\,
            I => \N__6251\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__6251\,
            I => \N__6245\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__6250\,
            I => \N__6241\
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__6249\,
            I => \N__6238\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__6248\,
            I => \N__6234\
        );

    \I__864\ : Span4Mux_h
    port map (
            O => \N__6245\,
            I => \N__6230\
        );

    \I__863\ : InMux
    port map (
            O => \N__6244\,
            I => \N__6217\
        );

    \I__862\ : InMux
    port map (
            O => \N__6241\,
            I => \N__6217\
        );

    \I__861\ : InMux
    port map (
            O => \N__6238\,
            I => \N__6217\
        );

    \I__860\ : InMux
    port map (
            O => \N__6237\,
            I => \N__6217\
        );

    \I__859\ : InMux
    port map (
            O => \N__6234\,
            I => \N__6217\
        );

    \I__858\ : InMux
    port map (
            O => \N__6233\,
            I => \N__6217\
        );

    \I__857\ : Odrv4
    port map (
            O => \N__6230\,
            I => \FSM_TEST_inst_RAPIDA.current_state_d_i_2\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__6217\,
            I => \FSM_TEST_inst_RAPIDA.current_state_d_i_2\
        );

    \I__855\ : InMux
    port map (
            O => \N__6212\,
            I => \N__6207\
        );

    \I__854\ : InMux
    port map (
            O => \N__6211\,
            I => \N__6204\
        );

    \I__853\ : InMux
    port map (
            O => \N__6210\,
            I => \N__6201\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__6207\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_7\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__6204\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_7\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__6201\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_7\
        );

    \I__849\ : CascadeMux
    port map (
            O => \N__6194\,
            I => \N__6191\
        );

    \I__848\ : InMux
    port map (
            O => \N__6191\,
            I => \N__6188\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__6188\,
            I => \FSM_TEST_inst_slow.flag_input_regZ0\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__6185\,
            I => \N__6181\
        );

    \I__845\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6177\
        );

    \I__844\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6174\
        );

    \I__843\ : InMux
    port map (
            O => \N__6180\,
            I => \N__6171\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__6177\,
            I => \N__6168\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__6174\,
            I => \N__6165\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__6171\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_6\
        );

    \I__839\ : Odrv4
    port map (
            O => \N__6168\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_6\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__6165\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_6\
        );

    \I__837\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6155\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__6155\,
            I => \FSM_TEST_inst_slow.current_state_RNO_3Z0Z_0\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__6152\,
            I => \FSM_TEST_inst_slow.current_state_RNO_4Z0Z_0_cascade_\
        );

    \I__834\ : InMux
    port map (
            O => \N__6149\,
            I => \N__6146\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__6146\,
            I => \FSM_TEST_inst_slow.current_state_RNO_5Z0Z_0\
        );

    \I__832\ : InMux
    port map (
            O => \N__6143\,
            I => \N__6140\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__6140\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_0\
        );

    \I__830\ : InMux
    port map (
            O => \N__6137\,
            I => \N__6134\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__6134\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_1\
        );

    \I__828\ : InMux
    port map (
            O => \N__6131\,
            I => \N__6128\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__6128\,
            I => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_2\
        );

    \I__826\ : InMux
    port map (
            O => \N__6125\,
            I => \N__6118\
        );

    \I__825\ : InMux
    port map (
            O => \N__6124\,
            I => \N__6118\
        );

    \I__824\ : InMux
    port map (
            O => \N__6123\,
            I => \N__6115\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__6118\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_0\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__6115\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_0\
        );

    \I__821\ : InMux
    port map (
            O => \N__6110\,
            I => \N__6107\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__6107\,
            I => \FSM_TEST_inst_slow.counter_stat_cry_1_THRU_CO\
        );

    \I__819\ : InMux
    port map (
            O => \N__6104\,
            I => \N__6097\
        );

    \I__818\ : InMux
    port map (
            O => \N__6103\,
            I => \N__6097\
        );

    \I__817\ : InMux
    port map (
            O => \N__6102\,
            I => \N__6094\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__6097\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_2\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__6094\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_2\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__6089\,
            I => \N__6086\
        );

    \I__813\ : InMux
    port map (
            O => \N__6086\,
            I => \N__6083\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__6083\,
            I => \FSM_TEST_inst_slow.counter_stat_cry_2_THRU_CO\
        );

    \I__811\ : InMux
    port map (
            O => \N__6080\,
            I => \N__6074\
        );

    \I__810\ : InMux
    port map (
            O => \N__6079\,
            I => \N__6069\
        );

    \I__809\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6069\
        );

    \I__808\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6066\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__6074\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_3\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__6069\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_3\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__6066\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_3\
        );

    \I__804\ : InMux
    port map (
            O => \N__6059\,
            I => \N__6056\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__6056\,
            I => \FSM_TEST_inst_slow.counter_stat_cry_0_THRU_CO\
        );

    \I__802\ : InMux
    port map (
            O => \N__6053\,
            I => \N__6048\
        );

    \I__801\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6045\
        );

    \I__800\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6042\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__6048\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_1\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__6045\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_1\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__6042\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_1\
        );

    \I__796\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6032\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__6032\,
            I => \FSM_TEST_inst_slow.counter_stat_cry_3_THRU_CO\
        );

    \I__794\ : InMux
    port map (
            O => \N__6029\,
            I => \N__6023\
        );

    \I__793\ : InMux
    port map (
            O => \N__6028\,
            I => \N__6020\
        );

    \I__792\ : InMux
    port map (
            O => \N__6027\,
            I => \N__6015\
        );

    \I__791\ : InMux
    port map (
            O => \N__6026\,
            I => \N__6015\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__6023\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_4\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__6020\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_4\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__6015\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_4\
        );

    \I__787\ : InMux
    port map (
            O => \N__6008\,
            I => \N__6002\
        );

    \I__786\ : InMux
    port map (
            O => \N__6007\,
            I => \N__5999\
        );

    \I__785\ : InMux
    port map (
            O => \N__6006\,
            I => \N__5994\
        );

    \I__784\ : InMux
    port map (
            O => \N__6005\,
            I => \N__5994\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__6002\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_4\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__5999\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_4\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5994\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_4\
        );

    \I__780\ : InMux
    port map (
            O => \N__5987\,
            I => \N__5981\
        );

    \I__779\ : InMux
    port map (
            O => \N__5986\,
            I => \N__5978\
        );

    \I__778\ : InMux
    port map (
            O => \N__5985\,
            I => \N__5975\
        );

    \I__777\ : InMux
    port map (
            O => \N__5984\,
            I => \N__5972\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__5981\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_5\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5978\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_5\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5975\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_5\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__5972\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_5\
        );

    \I__772\ : InMux
    port map (
            O => \N__5963\,
            I => \N__5959\
        );

    \I__771\ : InMux
    port map (
            O => \N__5962\,
            I => \N__5955\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5959\,
            I => \N__5952\
        );

    \I__769\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5949\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5955\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_1\
        );

    \I__767\ : Odrv4
    port map (
            O => \N__5952\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_1\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5949\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_1\
        );

    \I__765\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5939\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5939\,
            I => \N__5936\
        );

    \I__763\ : Odrv4
    port map (
            O => \N__5936\,
            I => \FSM_TEST_inst_RAPIDA.counter_idle_cry_0_THRU_CO\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__5933\,
            I => \FSM_TEST_inst_RAPIDA.N_126_1_i_cascade_\
        );

    \I__761\ : InMux
    port map (
            O => \N__5930\,
            I => \FSM_TEST_inst_slow.counter_stat_cry_0\
        );

    \I__760\ : InMux
    port map (
            O => \N__5927\,
            I => \FSM_TEST_inst_slow.counter_stat_cry_1\
        );

    \I__759\ : InMux
    port map (
            O => \N__5924\,
            I => \FSM_TEST_inst_slow.counter_stat_cry_2\
        );

    \I__758\ : InMux
    port map (
            O => \N__5921\,
            I => \FSM_TEST_inst_slow.counter_stat_cry_3\
        );

    \I__757\ : InMux
    port map (
            O => \N__5918\,
            I => \FSM_TEST_inst_slow.counter_stat_cry_4\
        );

    \I__756\ : InMux
    port map (
            O => \N__5915\,
            I => \FSM_TEST_inst_slow.counter_stat_cry_5\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__5912\,
            I => \N__5907\
        );

    \I__754\ : CascadeMux
    port map (
            O => \N__5911\,
            I => \N__5904\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__5910\,
            I => \N__5901\
        );

    \I__752\ : InMux
    port map (
            O => \N__5907\,
            I => \N__5898\
        );

    \I__751\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5895\
        );

    \I__750\ : InMux
    port map (
            O => \N__5901\,
            I => \N__5892\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__5898\,
            I => \N__5889\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5895\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_6\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__5892\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_6\
        );

    \I__746\ : Odrv4
    port map (
            O => \N__5889\,
            I => \FSM_TEST_inst_slow.counter_statZ0Z_6\
        );

    \I__745\ : CascadeMux
    port map (
            O => \N__5882\,
            I => \FSM_TEST_inst_slow.current_state_ns_0_a3_1_4_0_cascade_\
        );

    \I__744\ : InMux
    port map (
            O => \N__5879\,
            I => \N__5876\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__5876\,
            I => \FSM_TEST_inst_slow.current_state_ns_0_a3_1_5_0\
        );

    \I__742\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5870\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__5870\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_2\
        );

    \I__740\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5864\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__5864\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_3\
        );

    \I__738\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5858\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__5858\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_80\
        );

    \I__736\ : InMux
    port map (
            O => \N__5855\,
            I => \N__5852\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__5852\,
            I => \N__5849\
        );

    \I__734\ : Odrv4
    port map (
            O => \N__5849\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_42\
        );

    \I__733\ : InMux
    port map (
            O => \N__5846\,
            I => \N__5843\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__5843\,
            I => \N__5840\
        );

    \I__731\ : Odrv12
    port map (
            O => \N__5840\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_70\
        );

    \I__730\ : InMux
    port map (
            O => \N__5837\,
            I => \N__5834\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__5834\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_45\
        );

    \I__728\ : InMux
    port map (
            O => \N__5831\,
            I => \N__5828\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__5828\,
            I => \N__5825\
        );

    \I__726\ : Odrv4
    port map (
            O => \N__5825\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_76\
        );

    \I__725\ : InMux
    port map (
            O => \N__5822\,
            I => \N__5819\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5819\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_77\
        );

    \I__723\ : InMux
    port map (
            O => \N__5816\,
            I => \N__5813\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__5813\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_43\
        );

    \I__721\ : InMux
    port map (
            O => \N__5810\,
            I => \N__5807\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5807\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_44\
        );

    \I__719\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5801\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5801\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_78\
        );

    \I__717\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5795\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5795\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_79\
        );

    \I__715\ : InMux
    port map (
            O => \N__5792\,
            I => \N__5789\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__5789\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_13\
        );

    \I__713\ : InMux
    port map (
            O => \N__5786\,
            I => \N__5783\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__5783\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_0\
        );

    \I__711\ : InMux
    port map (
            O => \N__5780\,
            I => \N__5777\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5777\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_81\
        );

    \I__709\ : InMux
    port map (
            O => \N__5774\,
            I => \N__5771\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__5771\,
            I => \N__5768\
        );

    \I__707\ : Odrv4
    port map (
            O => \N__5768\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_46\
        );

    \I__706\ : InMux
    port map (
            O => \N__5765\,
            I => \N__5762\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__5762\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_4\
        );

    \I__704\ : InMux
    port map (
            O => \N__5759\,
            I => \N__5756\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__5756\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_1\
        );

    \I__702\ : CascadeMux
    port map (
            O => \N__5753\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2Z0Z_1_cascade_\
        );

    \I__701\ : InMux
    port map (
            O => \N__5750\,
            I => \N__5745\
        );

    \I__700\ : InMux
    port map (
            O => \N__5749\,
            I => \N__5742\
        );

    \I__699\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5739\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__5745\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_0\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5742\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_0\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5739\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_0\
        );

    \I__695\ : InMux
    port map (
            O => \N__5732\,
            I => \N__5729\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__5729\,
            I => \FSM_TEST_inst_RAPIDA.counter_stat_cry_0_THRU_CO\
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__5726\,
            I => \N__5721\
        );

    \I__692\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5715\
        );

    \I__691\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5704\
        );

    \I__690\ : InMux
    port map (
            O => \N__5721\,
            I => \N__5704\
        );

    \I__689\ : InMux
    port map (
            O => \N__5720\,
            I => \N__5704\
        );

    \I__688\ : InMux
    port map (
            O => \N__5719\,
            I => \N__5704\
        );

    \I__687\ : InMux
    port map (
            O => \N__5718\,
            I => \N__5704\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5715\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2Z0Z_1\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__5704\,
            I => \FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2Z0Z_1\
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__5699\,
            I => \N__5696\
        );

    \I__683\ : InMux
    port map (
            O => \N__5696\,
            I => \N__5693\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5693\,
            I => \FSM_TEST_inst_RAPIDA.counter_stat_cry_1_THRU_CO\
        );

    \I__681\ : InMux
    port map (
            O => \N__5690\,
            I => \N__5685\
        );

    \I__680\ : InMux
    port map (
            O => \N__5689\,
            I => \N__5682\
        );

    \I__679\ : InMux
    port map (
            O => \N__5688\,
            I => \N__5679\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__5685\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_2\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__5682\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_2\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__5679\,
            I => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_2\
        );

    \I__675\ : InMux
    port map (
            O => \N__5672\,
            I => \FSM_TEST_inst_RAPIDA.counter_idle_cry_0\
        );

    \I__674\ : InMux
    port map (
            O => \N__5669\,
            I => \FSM_TEST_inst_RAPIDA.counter_idle_cry_1\
        );

    \I__673\ : InMux
    port map (
            O => \N__5666\,
            I => \FSM_TEST_inst_RAPIDA.counter_idle_cry_2\
        );

    \I__672\ : InMux
    port map (
            O => \N__5663\,
            I => \FSM_TEST_inst_RAPIDA.counter_idle_cry_3\
        );

    \I__671\ : InMux
    port map (
            O => \N__5660\,
            I => \FSM_TEST_inst_RAPIDA.counter_idle_cry_4\
        );

    \I__670\ : InMux
    port map (
            O => \N__5657\,
            I => \N__5645\
        );

    \I__669\ : InMux
    port map (
            O => \N__5656\,
            I => \N__5645\
        );

    \I__668\ : InMux
    port map (
            O => \N__5655\,
            I => \N__5645\
        );

    \I__667\ : InMux
    port map (
            O => \N__5654\,
            I => \N__5645\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__5645\,
            I => \N__5638\
        );

    \I__665\ : InMux
    port map (
            O => \N__5644\,
            I => \N__5629\
        );

    \I__664\ : InMux
    port map (
            O => \N__5643\,
            I => \N__5629\
        );

    \I__663\ : InMux
    port map (
            O => \N__5642\,
            I => \N__5629\
        );

    \I__662\ : InMux
    port map (
            O => \N__5641\,
            I => \N__5629\
        );

    \I__661\ : Odrv4
    port map (
            O => \N__5638\,
            I => \FSM_TEST_inst_slow.N_134_1_i\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__5629\,
            I => \FSM_TEST_inst_slow.N_134_1_i\
        );

    \I__659\ : InMux
    port map (
            O => \N__5624\,
            I => \N__5619\
        );

    \I__658\ : InMux
    port map (
            O => \N__5623\,
            I => \N__5616\
        );

    \I__657\ : InMux
    port map (
            O => \N__5622\,
            I => \N__5613\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__5619\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_4\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__5616\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_4\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__5613\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_4\
        );

    \I__653\ : InMux
    port map (
            O => \N__5606\,
            I => \N__5601\
        );

    \I__652\ : InMux
    port map (
            O => \N__5605\,
            I => \N__5598\
        );

    \I__651\ : InMux
    port map (
            O => \N__5604\,
            I => \N__5595\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__5601\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_3\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__5598\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_3\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__5595\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_3\
        );

    \I__647\ : InMux
    port map (
            O => \N__5588\,
            I => \N__5585\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__5585\,
            I => \FSM_TEST_inst_RAPIDA.counter_stat_cry_3_THRU_CO\
        );

    \I__645\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__5579\,
            I => \FSM_TEST_inst_RAPIDA.counter_stat_cry_4_THRU_CO\
        );

    \I__643\ : InMux
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__5573\,
            I => \FSM_TEST_inst_RAPIDA.counter_stat_cry_2_THRU_CO\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__5570\,
            I => \FSM_TEST_inst_RAPIDA.counter_statlde_0_cascade_\
        );

    \I__640\ : InMux
    port map (
            O => \N__5567\,
            I => \FSM_TEST_inst_slow.counter_idle_cry_1\
        );

    \I__639\ : InMux
    port map (
            O => \N__5564\,
            I => \FSM_TEST_inst_slow.counter_idle_cry_2\
        );

    \I__638\ : InMux
    port map (
            O => \N__5561\,
            I => \FSM_TEST_inst_slow.counter_idle_cry_3\
        );

    \I__637\ : InMux
    port map (
            O => \N__5558\,
            I => \FSM_TEST_inst_slow.counter_idle_cry_4\
        );

    \I__636\ : InMux
    port map (
            O => \N__5555\,
            I => \FSM_TEST_inst_slow.counter_idle_cry_5\
        );

    \I__635\ : InMux
    port map (
            O => \N__5552\,
            I => \FSM_TEST_inst_slow.counter_idle_cry_6\
        );

    \I__634\ : CEMux
    port map (
            O => \N__5549\,
            I => \N__5546\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__5546\,
            I => \N__5543\
        );

    \I__632\ : Span4Mux_h
    port map (
            O => \N__5543\,
            I => \N__5540\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__5540\,
            I => \FSM_TEST_inst_slow.counter_idle_RNIHR3A2Z0Z_7\
        );

    \I__630\ : InMux
    port map (
            O => \N__5537\,
            I => \N__5533\
        );

    \I__629\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5530\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__5533\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_1\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__5530\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_1\
        );

    \I__626\ : InMux
    port map (
            O => \N__5525\,
            I => \N__5521\
        );

    \I__625\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5518\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__5521\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_2\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__5518\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_2\
        );

    \I__622\ : CascadeMux
    port map (
            O => \N__5513\,
            I => \N__5510\
        );

    \I__621\ : InMux
    port map (
            O => \N__5510\,
            I => \N__5506\
        );

    \I__620\ : InMux
    port map (
            O => \N__5509\,
            I => \N__5502\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__5506\,
            I => \N__5499\
        );

    \I__618\ : InMux
    port map (
            O => \N__5505\,
            I => \N__5496\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__5502\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_5\
        );

    \I__616\ : Odrv4
    port map (
            O => \N__5499\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_5\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__5496\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_5\
        );

    \I__614\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5485\
        );

    \I__613\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5482\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__5485\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_0\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__5482\,
            I => \FSM_TEST_inst_slow.counter_idleZ0Z_0\
        );

    \I__610\ : InMux
    port map (
            O => \N__5477\,
            I => \N__5474\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__5474\,
            I => \FSM_TEST_inst_slow.N_109_0\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__5471\,
            I => \N__5468\
        );

    \I__607\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5460\
        );

    \I__606\ : InMux
    port map (
            O => \N__5467\,
            I => \N__5460\
        );

    \I__605\ : InMux
    port map (
            O => \N__5466\,
            I => \N__5455\
        );

    \I__604\ : InMux
    port map (
            O => \N__5465\,
            I => \N__5455\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__5460\,
            I => \FSM_TEST_inst_slow.counter_dinZ0Z_0\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__5455\,
            I => \FSM_TEST_inst_slow.counter_dinZ0Z_0\
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__5450\,
            I => \N__5446\
        );

    \I__600\ : InMux
    port map (
            O => \N__5449\,
            I => \N__5442\
        );

    \I__599\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5437\
        );

    \I__598\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5437\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__5442\,
            I => \N__5432\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__5437\,
            I => \N__5432\
        );

    \I__595\ : Odrv4
    port map (
            O => \N__5432\,
            I => \FSM_TEST_inst_slow.counter_dinZ1Z_1\
        );

    \I__594\ : CascadeMux
    port map (
            O => \N__5429\,
            I => \FSM_TEST_inst_slow.N_134_1_cascade_\
        );

    \I__593\ : InMux
    port map (
            O => \N__5426\,
            I => \N__5423\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__5423\,
            I => \N__5420\
        );

    \I__591\ : Odrv4
    port map (
            O => \N__5420\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_15\
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__5417\,
            I => \N__5414\
        );

    \I__589\ : InMux
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__5411\,
            I => \N__5408\
        );

    \I__587\ : Span4Mux_v
    port map (
            O => \N__5408\,
            I => \N__5405\
        );

    \I__586\ : Odrv4
    port map (
            O => \N__5405\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_87\
        );

    \I__585\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5399\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__5399\,
            I => \FSM_TEST_inst_slow.G_31_1\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__5396\,
            I => \FSM_TEST_inst_slow.counter_statlde_0_cascade_\
        );

    \I__582\ : CEMux
    port map (
            O => \N__5393\,
            I => \N__5390\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__5390\,
            I => \N__5386\
        );

    \I__580\ : CEMux
    port map (
            O => \N__5389\,
            I => \N__5383\
        );

    \I__579\ : Span4Mux_h
    port map (
            O => \N__5386\,
            I => \N__5380\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__5383\,
            I => \N__5377\
        );

    \I__577\ : Span4Mux_h
    port map (
            O => \N__5380\,
            I => \N__5374\
        );

    \I__576\ : Odrv4
    port map (
            O => \N__5377\,
            I => \FSM_TEST_inst_slow.current_state_RNIR2L81Z0Z_1\
        );

    \I__575\ : Odrv4
    port map (
            O => \N__5374\,
            I => \FSM_TEST_inst_slow.current_state_RNIR2L81Z0Z_1\
        );

    \I__574\ : InMux
    port map (
            O => \N__5369\,
            I => \bfn_10_18_0_\
        );

    \I__573\ : InMux
    port map (
            O => \N__5366\,
            I => \FSM_TEST_inst_slow.counter_idle_cry_0\
        );

    \I__572\ : InMux
    port map (
            O => \N__5363\,
            I => \N__5360\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__5360\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_26\
        );

    \I__570\ : InMux
    port map (
            O => \N__5357\,
            I => \N__5354\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__5354\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_29\
        );

    \I__568\ : InMux
    port map (
            O => \N__5351\,
            I => \N__5348\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__5348\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_23\
        );

    \I__566\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5342\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__5342\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_24\
        );

    \I__564\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5336\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__5336\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_27\
        );

    \I__562\ : InMux
    port map (
            O => \N__5333\,
            I => \N__5330\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__5330\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_28\
        );

    \I__560\ : InMux
    port map (
            O => \N__5327\,
            I => \N__5324\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__5324\,
            I => \N__5321\
        );

    \I__558\ : Odrv4
    port map (
            O => \N__5321\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_47\
        );

    \I__557\ : InMux
    port map (
            O => \N__5318\,
            I => \N__5315\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__5315\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_73\
        );

    \I__555\ : InMux
    port map (
            O => \N__5312\,
            I => \N__5309\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__5309\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_74\
        );

    \I__553\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5303\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__5303\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_75\
        );

    \I__551\ : InMux
    port map (
            O => \N__5300\,
            I => \N__5297\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__5297\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_15\
        );

    \I__549\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5291\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__5291\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_14\
        );

    \I__547\ : InMux
    port map (
            O => \N__5288\,
            I => \N__5285\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__5285\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_22\
        );

    \I__545\ : InMux
    port map (
            O => \N__5282\,
            I => \N__5279\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__5279\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_20\
        );

    \I__543\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5273\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__5273\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_21\
        );

    \I__541\ : InMux
    port map (
            O => \N__5270\,
            I => \N__5267\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__5267\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_18\
        );

    \I__539\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5261\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__5261\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_19\
        );

    \I__537\ : InMux
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__5255\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_25\
        );

    \I__535\ : InMux
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__5249\,
            I => \FSM_TEST_inst_slow.CLK_uC_6jZ0Z_0\
        );

    \I__533\ : InMux
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__5243\,
            I => \N__5240\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__5240\,
            I => \FSM_TEST_inst_slow.CLK_uC_6gZ0Z_0\
        );

    \I__530\ : InMux
    port map (
            O => \N__5237\,
            I => \N__5234\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__5234\,
            I => \FSM_TEST_inst_slow.CLK_uC_6hZ0Z_0\
        );

    \I__528\ : InMux
    port map (
            O => \N__5231\,
            I => \FSM_TEST_inst_RAPIDA.counter_stat_cry_0\
        );

    \I__527\ : InMux
    port map (
            O => \N__5228\,
            I => \FSM_TEST_inst_RAPIDA.counter_stat_cry_1\
        );

    \I__526\ : InMux
    port map (
            O => \N__5225\,
            I => \FSM_TEST_inst_RAPIDA.counter_stat_cry_2\
        );

    \I__525\ : InMux
    port map (
            O => \N__5222\,
            I => \FSM_TEST_inst_RAPIDA.counter_stat_cry_3\
        );

    \I__524\ : InMux
    port map (
            O => \N__5219\,
            I => \FSM_TEST_inst_RAPIDA.counter_stat_cry_4\
        );

    \I__523\ : InMux
    port map (
            O => \N__5216\,
            I => \FSM_TEST_inst_RAPIDA.counter_stat_cry_5\
        );

    \I__522\ : InMux
    port map (
            O => \N__5213\,
            I => \N__5210\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__5210\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_7\
        );

    \I__520\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5204\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__5204\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_8\
        );

    \I__518\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5198\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__5198\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_9\
        );

    \I__516\ : InMux
    port map (
            O => \N__5195\,
            I => \N__5192\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__5192\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_10\
        );

    \I__514\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5186\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__5186\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_0\
        );

    \I__512\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5180\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__5180\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_1\
        );

    \I__510\ : InMux
    port map (
            O => \N__5177\,
            I => \N__5174\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__5174\,
            I => \FSM_TEST_inst_slow.CLK_uC_6iZ0Z_0\
        );

    \I__508\ : InMux
    port map (
            O => \N__5171\,
            I => \N__5168\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__5168\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_13\
        );

    \I__506\ : InMux
    port map (
            O => \N__5165\,
            I => \N__5162\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__5162\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_3\
        );

    \I__504\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5156\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__5156\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_2\
        );

    \I__502\ : InMux
    port map (
            O => \N__5153\,
            I => \N__5150\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__5150\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_11\
        );

    \I__500\ : InMux
    port map (
            O => \N__5147\,
            I => \N__5144\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__5144\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_14\
        );

    \I__498\ : InMux
    port map (
            O => \N__5141\,
            I => \N__5138\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__5138\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_4\
        );

    \I__496\ : InMux
    port map (
            O => \N__5135\,
            I => \N__5132\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__5132\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_5\
        );

    \I__494\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5126\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__5126\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_6\
        );

    \I__492\ : InMux
    port map (
            O => \N__5123\,
            I => \N__5120\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__5120\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_30\
        );

    \I__490\ : InMux
    port map (
            O => \N__5117\,
            I => \N__5114\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__5114\,
            I => \N__5111\
        );

    \I__488\ : Odrv4
    port map (
            O => \N__5111\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_71\
        );

    \I__487\ : InMux
    port map (
            O => \N__5108\,
            I => \N__5105\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__5105\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_31\
        );

    \I__485\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5099\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__5099\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_32\
        );

    \I__483\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5093\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__5093\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_72\
        );

    \I__481\ : InMux
    port map (
            O => \N__5090\,
            I => \N__5087\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__5087\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_41\
        );

    \I__479\ : InMux
    port map (
            O => \N__5084\,
            I => \N__5081\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__5081\,
            I => \N__5078\
        );

    \I__477\ : Span4Mux_v
    port map (
            O => \N__5078\,
            I => \N__5075\
        );

    \I__476\ : Odrv4
    port map (
            O => \N__5075\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_39\
        );

    \I__475\ : InMux
    port map (
            O => \N__5072\,
            I => \N__5069\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__5069\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_40\
        );

    \I__473\ : InMux
    port map (
            O => \N__5066\,
            I => \N__5063\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__5063\,
            I => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_12\
        );

    \I__471\ : InMux
    port map (
            O => \N__5060\,
            I => \N__5057\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__5057\,
            I => \FSM_TEST_inst_slow.CLK_uC_6eZ0Z_0\
        );

    \I__469\ : InMux
    port map (
            O => \N__5054\,
            I => \N__5051\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__5051\,
            I => \FSM_TEST_inst_slow.CLK_uC_6fZ0Z_0\
        );

    \I__467\ : InMux
    port map (
            O => \N__5048\,
            I => \N__5045\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__5045\,
            I => \FSM_TEST_inst_slow.CLK_uC_3_0_0\
        );

    \I__465\ : InMux
    port map (
            O => \N__5042\,
            I => \N__5039\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__5039\,
            I => \FSM_TEST_inst_slow.CLK_uC_4_0_0\
        );

    \I__463\ : InMux
    port map (
            O => \N__5036\,
            I => \N__5033\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__5033\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_16\
        );

    \I__461\ : InMux
    port map (
            O => \N__5030\,
            I => \N__5027\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__5027\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_17\
        );

    \I__459\ : InMux
    port map (
            O => \N__5024\,
            I => \N__5021\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__5021\,
            I => \N__5018\
        );

    \I__457\ : Odrv4
    port map (
            O => \N__5018\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_33\
        );

    \I__456\ : InMux
    port map (
            O => \N__5015\,
            I => \N__5012\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__5012\,
            I => \N__5009\
        );

    \I__454\ : Odrv4
    port map (
            O => \N__5009\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_48\
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__5006\,
            I => \N__5002\
        );

    \I__452\ : InMux
    port map (
            O => \N__5005\,
            I => \N__4997\
        );

    \I__451\ : InMux
    port map (
            O => \N__5002\,
            I => \N__4997\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4997\,
            I => \FSM_TEST_inst_slow.CLK_uCZ0\
        );

    \I__449\ : InMux
    port map (
            O => \N__4994\,
            I => \N__4991\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4991\,
            I => \FSM_TEST_inst_slow.CLK_uC_6c_0_0\
        );

    \I__447\ : InMux
    port map (
            O => \N__4988\,
            I => \N__4985\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__4985\,
            I => \FSM_TEST_inst_slow.CLK_uC_6b_0_0\
        );

    \I__445\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4979\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__4979\,
            I => \FSM_TEST_inst_slow.CLK_uC_2_0_0\
        );

    \I__443\ : InMux
    port map (
            O => \N__4976\,
            I => \N__4973\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4973\,
            I => \FSM_TEST_inst_slow.CLK_uC_5_0_0\
        );

    \I__441\ : InMux
    port map (
            O => \N__4970\,
            I => \N__4967\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4967\,
            I => \FSM_TEST_inst_slow.CLK_uC_6_0_0\
        );

    \I__439\ : InMux
    port map (
            O => \N__4964\,
            I => \N__4961\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__4961\,
            I => \FSM_TEST_inst_slow.CLK_uC_6dZ0Z_0\
        );

    \I__437\ : IoInMux
    port map (
            O => \N__4958\,
            I => \N__4955\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4955\,
            I => \N__4952\
        );

    \I__435\ : Span4Mux_s3_v
    port map (
            O => \N__4952\,
            I => \N__4949\
        );

    \I__434\ : Span4Mux_h
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__433\ : Odrv4
    port map (
            O => \N__4946\,
            I => \DYNCNF_i_0\
        );

    \I__432\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4940\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__4940\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_49\
        );

    \I__430\ : InMux
    port map (
            O => \N__4937\,
            I => \N__4934\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__4934\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_38\
        );

    \I__428\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4928\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__4928\,
            I => \N__4925\
        );

    \I__426\ : Odrv4
    port map (
            O => \N__4925\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_34\
        );

    \I__425\ : InMux
    port map (
            O => \N__4922\,
            I => \N__4919\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__4919\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_35\
        );

    \I__423\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4913\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__4913\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_36\
        );

    \I__421\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4907\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__4907\,
            I => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_37\
        );

    \I__419\ : IoInMux
    port map (
            O => \N__4904\,
            I => \N__4901\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__4901\,
            I => \N__4898\
        );

    \I__417\ : IoSpan4Mux
    port map (
            O => \N__4898\,
            I => \N__4895\
        );

    \I__416\ : Span4Mux_s3_v
    port map (
            O => \N__4895\,
            I => \N__4892\
        );

    \I__415\ : Sp12to4
    port map (
            O => \N__4892\,
            I => \N__4889\
        );

    \I__414\ : Span12Mux_v
    port map (
            O => \N__4889\,
            I => \N__4886\
        );

    \I__413\ : Span12Mux_v
    port map (
            O => \N__4886\,
            I => \N__4883\
        );

    \I__412\ : Odrv12
    port map (
            O => \N__4883\,
            I => \CLK_c\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_18_0_\
        );

    \RST_N_ibuf_RNIBJGC_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12008\,
            GLOBALBUFFEROUTPUT => \RST_N_c_i_g\
        );

    \FSM_TEST_inst_slow.current_state_RNIR2L81_1_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6737\,
            GLOBALBUFFEROUTPUT => \FSM_TEST_inst_slow.N_374_g\
        );

    \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIKIU51_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__11885\,
            GLOBALBUFFEROUTPUT => \FSM_TEST_inst_RAPIDA.N_256_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_36_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__7812\,
            in1 => \N__4922\,
            in2 => \_gnd_net_\,
            in3 => \N__8954\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10885\,
            ce => \N__7310\,
            sr => \N__10668\
        );

    \config_register_latched_dec_inst.DYNCNF_1_RNIP1121_0_0_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6791\,
            lcout => \DYNCNF_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_50_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__9049\,
            in1 => \_gnd_net_\,
            in2 => \N__7940\,
            in3 => \N__4943\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10868\,
            ce => \N__7313\,
            sr => \N__10671\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_49_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110100101"
        )
    port map (
            in0 => \N__9048\,
            in1 => \_gnd_net_\,
            in2 => \N__7939\,
            in3 => \N__5015\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10868\,
            ce => \N__7313\,
            sr => \N__10671\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_34_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5024\,
            in1 => \N__7931\,
            in2 => \_gnd_net_\,
            in3 => \N__9047\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10868\,
            ce => \N__7313\,
            sr => \N__10671\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_71_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__5846\,
            in1 => \N__7919\,
            in2 => \_gnd_net_\,
            in3 => \N__9046\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10874\,
            ce => \N__7312\,
            sr => \N__10669\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_39_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__4937\,
            in1 => \N__7887\,
            in2 => \_gnd_net_\,
            in3 => \N__8953\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10880\,
            ce => \N__7311\,
            sr => \N__10664\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_38_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__8952\,
            in1 => \N__4910\,
            in2 => \_gnd_net_\,
            in3 => \N__7888\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10880\,
            ce => \N__7311\,
            sr => \N__10664\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_35_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__4931\,
            in1 => \N__7885\,
            in2 => \_gnd_net_\,
            in3 => \N__8950\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10880\,
            ce => \N__7311\,
            sr => \N__10664\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_37_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__4916\,
            in1 => \N__7886\,
            in2 => \_gnd_net_\,
            in3 => \N__8951\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10880\,
            ce => \N__7311\,
            sr => \N__10664\
        );

    \FSM_TEST_inst_slow.CLK_uC_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011010010000"
        )
    port map (
            in0 => \N__7930\,
            in1 => \N__9045\,
            in2 => \N__5006\,
            in3 => \N__8546\,
            lcout => \FSM_TEST_inst_slow.CLK_uCZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10886\,
            ce => 'H',
            sr => \N__10659\
        );

    \FSM_TEST_inst_slow.CLK_uC_6d_0_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4994\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_6dZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10886\,
            ce => 'H',
            sr => \N__10659\
        );

    \FSM_TEST_inst_slow.CLK_uC_2_0_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5005\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10886\,
            ce => 'H',
            sr => \N__10659\
        );

    \FSM_TEST_inst_slow.CLK_uC_6c_0_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4988\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_6c_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10886\,
            ce => 'H',
            sr => \N__10659\
        );

    \FSM_TEST_inst_slow.CLK_uC_5_0_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5042\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10886\,
            ce => 'H',
            sr => \N__10659\
        );

    \FSM_TEST_inst_slow.CLK_uC_6b_0_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4970\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_6b_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10886\,
            ce => 'H',
            sr => \N__10659\
        );

    \FSM_TEST_inst_slow.CLK_uC_3_0_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4982\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10886\,
            ce => 'H',
            sr => \N__10659\
        );

    \FSM_TEST_inst_slow.CLK_uC_6_0_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4976\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10886\,
            ce => 'H',
            sr => \N__10659\
        );

    \FSM_TEST_inst_slow.CLK_uC_6e_0_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4964\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_6eZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10889\,
            ce => 'H',
            sr => \N__10654\
        );

    \FSM_TEST_inst_slow.CLK_uC_6f_0_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5060\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_6fZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10889\,
            ce => 'H',
            sr => \N__10654\
        );

    \FSM_TEST_inst_slow.CLK_uC_6g_0_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5054\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_6gZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10889\,
            ce => 'H',
            sr => \N__10654\
        );

    \FSM_TEST_inst_slow.CLK_uC_4_0_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5048\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10889\,
            ce => 'H',
            sr => \N__10654\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_16_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5300\,
            in1 => \N__7909\,
            in2 => \_gnd_net_\,
            in3 => \N__9060\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10839\,
            ce => \N__7323\,
            sr => \N__10672\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_17_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110100101"
        )
    port map (
            in0 => \N__9061\,
            in1 => \_gnd_net_\,
            in2 => \N__7938\,
            in3 => \N__5036\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10839\,
            ce => \N__7323\,
            sr => \N__10672\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_18_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__9041\,
            in1 => \N__5030\,
            in2 => \_gnd_net_\,
            in3 => \N__7848\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10847\,
            ce => \N__7319\,
            sr => \N__10670\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_33_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5102\,
            in1 => \N__7841\,
            in2 => \_gnd_net_\,
            in3 => \N__9027\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10855\,
            ce => \N__7316\,
            sr => \N__10665\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_41_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__9028\,
            in1 => \_gnd_net_\,
            in2 => \N__7921\,
            in3 => \N__5072\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10855\,
            ce => \N__7316\,
            sr => \N__10665\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_31_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110100101"
        )
    port map (
            in0 => \N__9026\,
            in1 => \_gnd_net_\,
            in2 => \N__7920\,
            in3 => \N__5123\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10855\,
            ce => \N__7316\,
            sr => \N__10665\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_48_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__9029\,
            in1 => \_gnd_net_\,
            in2 => \N__7922\,
            in3 => \N__5327\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10855\,
            ce => \N__7316\,
            sr => \N__10665\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_30_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5357\,
            in1 => \N__7837\,
            in2 => \_gnd_net_\,
            in3 => \N__9025\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10855\,
            ce => \N__7316\,
            sr => \N__10665\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_72_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__8987\,
            in1 => \_gnd_net_\,
            in2 => \N__7917\,
            in3 => \N__5117\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10862\,
            ce => \N__7314\,
            sr => \N__10660\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_32_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__5108\,
            in1 => \N__8984\,
            in2 => \_gnd_net_\,
            in3 => \N__7813\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10862\,
            ce => \N__7314\,
            sr => \N__10660\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_73_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__8988\,
            in1 => \_gnd_net_\,
            in2 => \N__7918\,
            in3 => \N__5096\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10862\,
            ce => \N__7314\,
            sr => \N__10660\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_42_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110100101"
        )
    port map (
            in0 => \N__8986\,
            in1 => \_gnd_net_\,
            in2 => \N__7916\,
            in3 => \N__5090\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10862\,
            ce => \N__7314\,
            sr => \N__10660\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_40_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__5084\,
            in1 => \N__8985\,
            in2 => \_gnd_net_\,
            in3 => \N__7814\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10862\,
            ce => \N__7314\,
            sr => \N__10660\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_13_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__7665\,
            in1 => \N__5066\,
            in2 => \_gnd_net_\,
            in3 => \N__8932\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10869\,
            ce => \N__5393\,
            sr => \N__10655\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_4_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__8937\,
            in1 => \N__5165\,
            in2 => \_gnd_net_\,
            in3 => \N__7670\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10869\,
            ce => \N__5393\,
            sr => \N__10655\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_12_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__7664\,
            in1 => \N__5153\,
            in2 => \_gnd_net_\,
            in3 => \N__8931\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10869\,
            ce => \N__5393\,
            sr => \N__10655\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_14_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__8933\,
            in1 => \N__5171\,
            in2 => \_gnd_net_\,
            in3 => \N__7666\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10869\,
            ce => \N__5393\,
            sr => \N__10655\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_3_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__7669\,
            in1 => \N__5159\,
            in2 => \_gnd_net_\,
            in3 => \N__8936\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10869\,
            ce => \N__5393\,
            sr => \N__10655\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_2_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__8935\,
            in1 => \N__5183\,
            in2 => \_gnd_net_\,
            in3 => \N__7668\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10869\,
            ce => \N__5393\,
            sr => \N__10655\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_11_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__7663\,
            in1 => \N__5195\,
            in2 => \_gnd_net_\,
            in3 => \N__8930\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10869\,
            ce => \N__5393\,
            sr => \N__10655\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_15_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__8934\,
            in1 => \N__5147\,
            in2 => \_gnd_net_\,
            in3 => \N__7667\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10869\,
            ce => \N__5393\,
            sr => \N__10655\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_6_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__9008\,
            in1 => \N__5135\,
            in2 => \_gnd_net_\,
            in3 => \N__7834\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10875\,
            ce => \N__5389\,
            sr => \N__10650\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_5_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__5141\,
            in1 => \N__7831\,
            in2 => \_gnd_net_\,
            in3 => \N__9007\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10875\,
            ce => \N__5389\,
            sr => \N__10650\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_7_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__9009\,
            in1 => \N__5129\,
            in2 => \_gnd_net_\,
            in3 => \N__7835\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10875\,
            ce => \N__5389\,
            sr => \N__10650\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_0_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7829\,
            in2 => \_gnd_net_\,
            in3 => \N__9004\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10875\,
            ce => \N__5389\,
            sr => \N__10650\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_8_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__9010\,
            in1 => \N__5213\,
            in2 => \_gnd_net_\,
            in3 => \N__7836\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10875\,
            ce => \N__5389\,
            sr => \N__10650\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_9_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5207\,
            in1 => \N__7832\,
            in2 => \_gnd_net_\,
            in3 => \N__9011\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10875\,
            ce => \N__5389\,
            sr => \N__10650\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_10_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__9005\,
            in1 => \N__5201\,
            in2 => \_gnd_net_\,
            in3 => \N__7833\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10875\,
            ce => \N__5389\,
            sr => \N__10650\
        );

    \FSM_TEST_inst_slow.bit_sequence_din_1_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__5189\,
            in1 => \N__7830\,
            in2 => \_gnd_net_\,
            in3 => \N__9006\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10875\,
            ce => \N__5389\,
            sr => \N__10650\
        );

    \FSM_TEST_inst_slow.counter_din_1_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110110000000"
        )
    port map (
            in0 => \N__7239\,
            in1 => \N__6718\,
            in2 => \N__5471\,
            in3 => \N__5449\,
            lcout => \FSM_TEST_inst_slow.counter_dinZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10881\,
            ce => 'H',
            sr => \N__10646\
        );

    \FSM_TEST_inst_slow.counter_din_0_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011001100"
        )
    port map (
            in0 => \N__6717\,
            in1 => \N__5467\,
            in2 => \_gnd_net_\,
            in3 => \N__7238\,
            lcout => \FSM_TEST_inst_slow.counter_dinZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10881\,
            ce => 'H',
            sr => \N__10646\
        );

    \FSM_TEST_inst_slow.counter_din_3_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101100011010000"
        )
    port map (
            in0 => \N__7240\,
            in1 => \N__6719\,
            in2 => \N__6942\,
            in3 => \N__5477\,
            lcout => \FSM_TEST_inst_slow.counter_dinZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10881\,
            ce => 'H',
            sr => \N__10646\
        );

    \FSM_TEST_inst_slow.CLK_uC_6i_0_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5237\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_6iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10881\,
            ce => 'H',
            sr => \N__10646\
        );

    \FSM_TEST_inst_slow.CLK_uC_6j_0_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5177\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_6jZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10881\,
            ce => 'H',
            sr => \N__10646\
        );

    \FSM_TEST_inst_slow.CLK_uC_6k_0_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5252\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_6kZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10881\,
            ce => 'H',
            sr => \N__10646\
        );

    \FSM_TEST_inst_slow.CLK_uC_6h_0_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5246\,
            lcout => \FSM_TEST_inst_slow.CLK_uC_6hZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10881\,
            ce => 'H',
            sr => \N__10646\
        );

    \FSM_TEST_inst_RAPIDA.counter_stat_cry_c_0_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5748\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \FSM_TEST_inst_RAPIDA.counter_stat_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_stat_cry_0_THRU_LUT4_0_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5958\,
            in2 => \_gnd_net_\,
            in3 => \N__5231\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_stat_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_RAPIDA.counter_stat_cry_0\,
            carryout => \FSM_TEST_inst_RAPIDA.counter_stat_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_stat_cry_1_THRU_LUT4_0_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5688\,
            in2 => \_gnd_net_\,
            in3 => \N__5228\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_stat_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_RAPIDA.counter_stat_cry_1\,
            carryout => \FSM_TEST_inst_RAPIDA.counter_stat_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_stat_cry_2_THRU_LUT4_0_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6985\,
            in2 => \_gnd_net_\,
            in3 => \N__5225\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_stat_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_RAPIDA.counter_stat_cry_2\,
            carryout => \FSM_TEST_inst_RAPIDA.counter_stat_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_stat_cry_3_THRU_LUT4_0_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6007\,
            in2 => \_gnd_net_\,
            in3 => \N__5222\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_stat_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_RAPIDA.counter_stat_cry_3\,
            carryout => \FSM_TEST_inst_RAPIDA.counter_stat_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_stat_cry_4_THRU_LUT4_0_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5986\,
            in2 => \_gnd_net_\,
            in3 => \N__5219\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_stat_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_RAPIDA.counter_stat_cry_4\,
            carryout => \FSM_TEST_inst_RAPIDA.counter_stat_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_stat_6_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011010001110000"
        )
    port map (
            in0 => \N__6254\,
            in1 => \N__5725\,
            in2 => \N__7021\,
            in3 => \N__5216\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10887\,
            ce => 'H',
            sr => \N__10641\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_87_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__6578\,
            in1 => \N__7929\,
            in2 => \_gnd_net_\,
            in3 => \N__9062\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10821\,
            ce => \N__7331\,
            sr => \N__10673\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_15_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__5294\,
            in1 => \N__7908\,
            in2 => \_gnd_net_\,
            in3 => \N__9051\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10826\,
            ce => \N__7324\,
            sr => \N__10666\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_14_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5792\,
            in1 => \N__7907\,
            in2 => \_gnd_net_\,
            in3 => \N__9050\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10826\,
            ce => \N__7324\,
            sr => \N__10666\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_23_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__9024\,
            in1 => \N__5288\,
            in2 => \_gnd_net_\,
            in3 => \N__7881\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10832\,
            ce => \N__7320\,
            sr => \N__10661\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_20_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__7878\,
            in1 => \N__5264\,
            in2 => \_gnd_net_\,
            in3 => \N__9021\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10832\,
            ce => \N__7320\,
            sr => \N__10661\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_22_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__7880\,
            in1 => \N__5276\,
            in2 => \_gnd_net_\,
            in3 => \N__9023\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10832\,
            ce => \N__7320\,
            sr => \N__10661\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_21_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__9022\,
            in1 => \N__5282\,
            in2 => \_gnd_net_\,
            in3 => \N__7879\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10832\,
            ce => \N__7320\,
            sr => \N__10661\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_19_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__7877\,
            in1 => \N__5270\,
            in2 => \_gnd_net_\,
            in3 => \N__9020\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10832\,
            ce => \N__7320\,
            sr => \N__10661\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_26_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__9015\,
            in1 => \_gnd_net_\,
            in2 => \N__7926\,
            in3 => \N__5258\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10841\,
            ce => \N__7317\,
            sr => \N__10656\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_25_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__5345\,
            in1 => \N__7865\,
            in2 => \_gnd_net_\,
            in3 => \N__9014\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10841\,
            ce => \N__7317\,
            sr => \N__10656\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_27_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__9016\,
            in1 => \_gnd_net_\,
            in2 => \N__7927\,
            in3 => \N__5363\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10841\,
            ce => \N__7317\,
            sr => \N__10656\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_29_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5333\,
            in1 => \N__7875\,
            in2 => \_gnd_net_\,
            in3 => \N__9018\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10841\,
            ce => \N__7317\,
            sr => \N__10656\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_24_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5351\,
            in1 => \N__7864\,
            in2 => \_gnd_net_\,
            in3 => \N__9013\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10841\,
            ce => \N__7317\,
            sr => \N__10656\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_28_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110100101"
        )
    port map (
            in0 => \N__9017\,
            in1 => \_gnd_net_\,
            in2 => \N__7928\,
            in3 => \N__5339\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10841\,
            ce => \N__7317\,
            sr => \N__10656\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_47_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5774\,
            in1 => \N__7876\,
            in2 => \_gnd_net_\,
            in3 => \N__9019\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10841\,
            ce => \N__7317\,
            sr => \N__10656\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_76_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5306\,
            in1 => \N__7863\,
            in2 => \_gnd_net_\,
            in3 => \N__8983\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10849\,
            ce => \N__7315\,
            sr => \N__10651\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_74_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5318\,
            in1 => \N__7859\,
            in2 => \_gnd_net_\,
            in3 => \N__8981\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10849\,
            ce => \N__7315\,
            sr => \N__10651\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_75_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__8982\,
            in1 => \_gnd_net_\,
            in2 => \N__7925\,
            in3 => \N__5312\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10849\,
            ce => \N__7315\,
            sr => \N__10651\
        );

    \FSM_TEST_inst_slow.current_state_RNIV6JP_2_1_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7639\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8854\,
            lcout => OPEN,
            ltout => \FSM_TEST_inst_slow.N_134_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.counter_idle_RNIHR3A2_7_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100000000"
        )
    port map (
            in0 => \N__6211\,
            in1 => \N__5402\,
            in2 => \N__5429\,
            in3 => \N__7227\,
            lcout => \FSM_TEST_inst_slow.counter_idle_RNIHR3A2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.MOSI_er_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__7644\,
            in1 => \N__5426\,
            in2 => \N__5417\,
            in3 => \N__8857\,
            lcout => mosi_slow,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10856\,
            ce => \N__7241\,
            sr => \N__10647\
        );

    \FSM_TEST_inst_slow.counter_idle_RNIMHOQ_3_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011111"
        )
    port map (
            in0 => \N__5605\,
            in1 => \N__5623\,
            in2 => \N__6185\,
            in3 => \N__5505\,
            lcout => \FSM_TEST_inst_slow.G_31_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.counter_stat_RNIE9EB1_6_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__9192\,
            in1 => \N__6026\,
            in2 => \N__5912\,
            in3 => \N__6077\,
            lcout => OPEN,
            ltout => \FSM_TEST_inst_slow.counter_statlde_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.current_state_RNI9C3K2_1_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100000000"
        )
    port map (
            in0 => \N__8855\,
            in1 => \N__7640\,
            in2 => \N__5396\,
            in3 => \N__7225\,
            lcout => \FSM_TEST_inst_slow.current_state_RNI9C3K2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.current_state_RNIR2L81_1_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001010"
        )
    port map (
            in0 => \N__7226\,
            in1 => \_gnd_net_\,
            in2 => \N__7828\,
            in3 => \N__8856\,
            lcout => \FSM_TEST_inst_slow.current_state_RNIR2L81Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.current_state_RNO_7_0_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6027\,
            in1 => \N__6052\,
            in2 => \N__9197\,
            in3 => \N__7638\,
            lcout => \FSM_TEST_inst_slow.current_state_ns_0_a3_1_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.counter_idle_0_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5654\,
            in1 => \N__5489\,
            in2 => \_gnd_net_\,
            in3 => \N__5369\,
            lcout => \FSM_TEST_inst_slow.counter_idleZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_18_0_\,
            carryout => \FSM_TEST_inst_slow.counter_idle_cry_0\,
            clk => \N__10863\,
            ce => \N__5549\,
            sr => \N__10642\
        );

    \FSM_TEST_inst_slow.counter_idle_1_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5641\,
            in1 => \N__5537\,
            in2 => \_gnd_net_\,
            in3 => \N__5366\,
            lcout => \FSM_TEST_inst_slow.counter_idleZ0Z_1\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_slow.counter_idle_cry_0\,
            carryout => \FSM_TEST_inst_slow.counter_idle_cry_1\,
            clk => \N__10863\,
            ce => \N__5549\,
            sr => \N__10642\
        );

    \FSM_TEST_inst_slow.counter_idle_2_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5655\,
            in1 => \N__5525\,
            in2 => \_gnd_net_\,
            in3 => \N__5567\,
            lcout => \FSM_TEST_inst_slow.counter_idleZ0Z_2\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_slow.counter_idle_cry_1\,
            carryout => \FSM_TEST_inst_slow.counter_idle_cry_2\,
            clk => \N__10863\,
            ce => \N__5549\,
            sr => \N__10642\
        );

    \FSM_TEST_inst_slow.counter_idle_3_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5642\,
            in1 => \N__5606\,
            in2 => \_gnd_net_\,
            in3 => \N__5564\,
            lcout => \FSM_TEST_inst_slow.counter_idleZ0Z_3\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_slow.counter_idle_cry_2\,
            carryout => \FSM_TEST_inst_slow.counter_idle_cry_3\,
            clk => \N__10863\,
            ce => \N__5549\,
            sr => \N__10642\
        );

    \FSM_TEST_inst_slow.counter_idle_4_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5656\,
            in1 => \N__5624\,
            in2 => \_gnd_net_\,
            in3 => \N__5561\,
            lcout => \FSM_TEST_inst_slow.counter_idleZ0Z_4\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_slow.counter_idle_cry_3\,
            carryout => \FSM_TEST_inst_slow.counter_idle_cry_4\,
            clk => \N__10863\,
            ce => \N__5549\,
            sr => \N__10642\
        );

    \FSM_TEST_inst_slow.counter_idle_5_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5643\,
            in1 => \N__5509\,
            in2 => \_gnd_net_\,
            in3 => \N__5558\,
            lcout => \FSM_TEST_inst_slow.counter_idleZ0Z_5\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_slow.counter_idle_cry_4\,
            carryout => \FSM_TEST_inst_slow.counter_idle_cry_5\,
            clk => \N__10863\,
            ce => \N__5549\,
            sr => \N__10642\
        );

    \FSM_TEST_inst_slow.counter_idle_6_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5657\,
            in1 => \N__6180\,
            in2 => \_gnd_net_\,
            in3 => \N__5555\,
            lcout => \FSM_TEST_inst_slow.counter_idleZ0Z_6\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_slow.counter_idle_cry_5\,
            carryout => \FSM_TEST_inst_slow.counter_idle_cry_6\,
            clk => \N__10863\,
            ce => \N__5549\,
            sr => \N__10642\
        );

    \FSM_TEST_inst_slow.counter_idle_7_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5644\,
            in1 => \N__6212\,
            in2 => \_gnd_net_\,
            in3 => \N__5552\,
            lcout => \FSM_TEST_inst_slow.counter_idleZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10863\,
            ce => \N__5549\,
            sr => \N__10642\
        );

    \FSM_TEST_inst_slow.current_state_RNO_3_0_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__5536\,
            in1 => \N__5524\,
            in2 => \N__5513\,
            in3 => \N__5488\,
            lcout => \FSM_TEST_inst_slow.current_state_RNO_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.counter_din_RNO_0_3_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__5466\,
            in1 => \_gnd_net_\,
            in2 => \N__5450\,
            in3 => \N__6920\,
            lcout => \FSM_TEST_inst_slow.N_109_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.counter_din_RNID6M9_1_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5465\,
            in2 => \_gnd_net_\,
            in3 => \N__5445\,
            lcout => \FSM_TEST_inst_slow.N_106_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.current_state_RNO_4_0_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5689\,
            in2 => \_gnd_net_\,
            in3 => \N__5749\,
            lcout => \FSM_TEST_inst_RAPIDA.G_24_0_a4_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.current_state_RNIV6JP_0_1_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9003\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7850\,
            lcout => \FSM_TEST_inst_slow.current_state_d_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.current_state_RNIV6JP_1_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7849\,
            in2 => \_gnd_net_\,
            in3 => \N__9002\,
            lcout => \FSM_TEST_inst_slow.N_134_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.current_state_RNO_5_0_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5622\,
            in2 => \_gnd_net_\,
            in3 => \N__5604\,
            lcout => \FSM_TEST_inst_slow.current_state_RNO_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_stat_4_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010011000101010"
        )
    port map (
            in0 => \N__6006\,
            in1 => \N__5720\,
            in2 => \N__6250\,
            in3 => \N__5588\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10876\,
            ce => 'H',
            sr => \N__10634\
        );

    \FSM_TEST_inst_RAPIDA.counter_stat_5_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001111100100000"
        )
    port map (
            in0 => \N__5582\,
            in1 => \N__6244\,
            in2 => \N__5726\,
            in3 => \N__5987\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10876\,
            ce => 'H',
            sr => \N__10634\
        );

    \FSM_TEST_inst_RAPIDA.counter_stat_3_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011010101010"
        )
    port map (
            in0 => \N__6984\,
            in1 => \N__5576\,
            in2 => \N__6249\,
            in3 => \N__5724\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10876\,
            ce => 'H',
            sr => \N__10634\
        );

    \FSM_TEST_inst_RAPIDA.counter_stat_RNIUUIP1_6_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__5984\,
            in1 => \N__6005\,
            in2 => \N__7017\,
            in3 => \N__6983\,
            lcout => OPEN,
            ltout => \FSM_TEST_inst_RAPIDA.counter_statlde_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2_1_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001001100"
        )
    port map (
            in0 => \N__9412\,
            in1 => \N__11649\,
            in2 => \N__5570\,
            in3 => \N__11459\,
            lcout => \FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2Z0Z_1\,
            ltout => \FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_stat_0_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001111100100000"
        )
    port map (
            in0 => \N__6616\,
            in1 => \N__6233\,
            in2 => \N__5753\,
            in3 => \N__5750\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10876\,
            ce => 'H',
            sr => \N__10634\
        );

    \FSM_TEST_inst_RAPIDA.counter_stat_1_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011011100001000"
        )
    port map (
            in0 => \N__5732\,
            in1 => \N__5719\,
            in2 => \N__6248\,
            in3 => \N__5962\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10876\,
            ce => 'H',
            sr => \N__10634\
        );

    \FSM_TEST_inst_RAPIDA.counter_stat_2_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101011100100000"
        )
    port map (
            in0 => \N__5718\,
            in1 => \N__6237\,
            in2 => \N__5699\,
            in3 => \N__5690\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_statZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10876\,
            ce => 'H',
            sr => \N__10634\
        );

    \FSM_TEST_inst_RAPIDA.counter_idle_cry_c_0_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6417\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => \FSM_TEST_inst_RAPIDA.counter_idle_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_idle_cry_0_THRU_LUT4_0_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6460\,
            in2 => \_gnd_net_\,
            in3 => \N__5672\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_idle_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_RAPIDA.counter_idle_cry_0\,
            carryout => \FSM_TEST_inst_RAPIDA.counter_idle_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_idle_cry_1_THRU_LUT4_0_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6439\,
            in2 => \_gnd_net_\,
            in3 => \N__5669\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_idle_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_RAPIDA.counter_idle_cry_1\,
            carryout => \FSM_TEST_inst_RAPIDA.counter_idle_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_idle_cry_2_THRU_LUT4_0_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6298\,
            in2 => \_gnd_net_\,
            in3 => \N__5666\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_idle_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_RAPIDA.counter_idle_cry_2\,
            carryout => \FSM_TEST_inst_RAPIDA.counter_idle_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_idle_cry_3_THRU_LUT4_0_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6317\,
            in2 => \_gnd_net_\,
            in3 => \N__5663\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_idle_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_RAPIDA.counter_idle_cry_3\,
            carryout => \FSM_TEST_inst_RAPIDA.counter_idle_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_idle_5_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001110001001100"
        )
    port map (
            in0 => \N__6484\,
            in1 => \N__6276\,
            in2 => \N__6528\,
            in3 => \N__5660\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10882\,
            ce => 'H',
            sr => \N__10629\
        );

    \FSM_TEST_inst_RAPIDA.flag_input_reg_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6602\,
            lcout => \FSM_TEST_inst_RAPIDA.flag_input_regZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10888\,
            ce => 'H',
            sr => \N__10624\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_13_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__8980\,
            in1 => \N__6545\,
            in2 => \_gnd_net_\,
            in3 => \N__7827\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10823\,
            ce => \N__7328\,
            sr => \N__10662\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_1_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110100101"
        )
    port map (
            in0 => \N__8956\,
            in1 => \_gnd_net_\,
            in2 => \N__7923\,
            in3 => \N__5786\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10827\,
            ce => \N__7325\,
            sr => \N__10657\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_82_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__5780\,
            in1 => \N__7858\,
            in2 => \_gnd_net_\,
            in3 => \N__8958\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10827\,
            ce => \N__7325\,
            sr => \N__10657\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_0_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7851\,
            in2 => \_gnd_net_\,
            in3 => \N__8955\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10827\,
            ce => \N__7325\,
            sr => \N__10657\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_81_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110100101"
        )
    port map (
            in0 => \N__8957\,
            in1 => \_gnd_net_\,
            in2 => \N__7924\,
            in3 => \N__5861\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10827\,
            ce => \N__7325\,
            sr => \N__10657\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_46_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__8973\,
            in1 => \_gnd_net_\,
            in2 => \N__7901\,
            in3 => \N__5837\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10833\,
            ce => \N__7321\,
            sr => \N__10652\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_4_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__5867\,
            in1 => \N__7766\,
            in2 => \_gnd_net_\,
            in3 => \N__8974\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10833\,
            ce => \N__7321\,
            sr => \N__10652\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_5_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110100101"
        )
    port map (
            in0 => \N__8975\,
            in1 => \_gnd_net_\,
            in2 => \N__7902\,
            in3 => \N__5765\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10833\,
            ce => \N__7321\,
            sr => \N__10652\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_2_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5759\,
            in1 => \N__7761\,
            in2 => \_gnd_net_\,
            in3 => \N__8971\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10833\,
            ce => \N__7321\,
            sr => \N__10652\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_3_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__5873\,
            in1 => \N__7762\,
            in2 => \_gnd_net_\,
            in3 => \N__8972\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10833\,
            ce => \N__7321\,
            sr => \N__10652\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_80_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__8976\,
            in1 => \_gnd_net_\,
            in2 => \N__7903\,
            in3 => \N__5798\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10833\,
            ce => \N__7321\,
            sr => \N__10652\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_43_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5855\,
            in1 => \N__7561\,
            in2 => \_gnd_net_\,
            in3 => \N__8713\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10842\,
            ce => \N__7318\,
            sr => \N__10648\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_70_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__6758\,
            in1 => \N__7563\,
            in2 => \_gnd_net_\,
            in3 => \N__8716\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10842\,
            ce => \N__7318\,
            sr => \N__10648\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_45_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__8715\,
            in1 => \N__5810\,
            in2 => \_gnd_net_\,
            in3 => \N__7565\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10842\,
            ce => \N__7318\,
            sr => \N__10648\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_77_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5831\,
            in1 => \N__7564\,
            in2 => \_gnd_net_\,
            in3 => \N__8717\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10842\,
            ce => \N__7318\,
            sr => \N__10648\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_78_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__8718\,
            in1 => \N__5822\,
            in2 => \_gnd_net_\,
            in3 => \N__7566\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10842\,
            ce => \N__7318\,
            sr => \N__10648\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_44_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__5816\,
            in1 => \N__7562\,
            in2 => \_gnd_net_\,
            in3 => \N__8714\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10842\,
            ce => \N__7318\,
            sr => \N__10648\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_79_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__8719\,
            in1 => \N__5804\,
            in2 => \_gnd_net_\,
            in3 => \N__7567\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10842\,
            ce => \N__7318\,
            sr => \N__10648\
        );

    \FSM_TEST_inst_slow.counter_stat_cry_c_0_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6123\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \FSM_TEST_inst_slow.counter_stat_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.counter_stat_cry_0_THRU_LUT4_0_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6051\,
            in2 => \_gnd_net_\,
            in3 => \N__5930\,
            lcout => \FSM_TEST_inst_slow.counter_stat_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_slow.counter_stat_cry_0\,
            carryout => \FSM_TEST_inst_slow.counter_stat_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.counter_stat_cry_1_THRU_LUT4_0_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6102\,
            in2 => \_gnd_net_\,
            in3 => \N__5927\,
            lcout => \FSM_TEST_inst_slow.counter_stat_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_slow.counter_stat_cry_1\,
            carryout => \FSM_TEST_inst_slow.counter_stat_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.counter_stat_cry_2_THRU_LUT4_0_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6080\,
            in2 => \_gnd_net_\,
            in3 => \N__5924\,
            lcout => \FSM_TEST_inst_slow.counter_stat_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_slow.counter_stat_cry_2\,
            carryout => \FSM_TEST_inst_slow.counter_stat_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.counter_stat_cry_3_THRU_LUT4_0_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6028\,
            in2 => \_gnd_net_\,
            in3 => \N__5921\,
            lcout => \FSM_TEST_inst_slow.counter_stat_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_slow.counter_stat_cry_3\,
            carryout => \FSM_TEST_inst_slow.counter_stat_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.counter_stat_cry_4_THRU_LUT4_0_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9196\,
            in2 => \_gnd_net_\,
            in3 => \N__5918\,
            lcout => \FSM_TEST_inst_slow.counter_stat_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \FSM_TEST_inst_slow.counter_stat_cry_4\,
            carryout => \FSM_TEST_inst_slow.counter_stat_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.counter_stat_6_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011010001110000"
        )
    port map (
            in0 => \N__9250\,
            in1 => \N__9293\,
            in2 => \N__5911\,
            in3 => \N__5915\,
            lcout => \FSM_TEST_inst_slow.counter_statZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10850\,
            ce => 'H',
            sr => \N__10643\
        );

    \FSM_TEST_inst_slow.current_state_RNO_6_0_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6103\,
            in1 => \N__6078\,
            in2 => \N__5910\,
            in3 => \N__6124\,
            lcout => OPEN,
            ltout => \FSM_TEST_inst_slow.current_state_ns_0_a3_1_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.current_state_RNO_1_0_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5882\,
            in3 => \N__5879\,
            lcout => \FSM_TEST_inst_slow.current_state_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.counter_stat_0_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101011100100000"
        )
    port map (
            in0 => \N__9287\,
            in1 => \N__9239\,
            in2 => \N__6617\,
            in3 => \N__6125\,
            lcout => \FSM_TEST_inst_slow.counter_statZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10857\,
            ce => 'H',
            sr => \N__10638\
        );

    \FSM_TEST_inst_slow.counter_stat_2_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011011001100"
        )
    port map (
            in0 => \N__6110\,
            in1 => \N__6104\,
            in2 => \N__9255\,
            in3 => \N__9291\,
            lcout => \FSM_TEST_inst_slow.counter_statZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10857\,
            ce => 'H',
            sr => \N__10638\
        );

    \FSM_TEST_inst_slow.counter_stat_3_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101011100100000"
        )
    port map (
            in0 => \N__9288\,
            in1 => \N__9240\,
            in2 => \N__6089\,
            in3 => \N__6079\,
            lcout => \FSM_TEST_inst_slow.counter_statZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10857\,
            ce => 'H',
            sr => \N__10638\
        );

    \FSM_TEST_inst_slow.counter_stat_1_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011011100001000"
        )
    port map (
            in0 => \N__6059\,
            in1 => \N__9290\,
            in2 => \N__9254\,
            in3 => \N__6053\,
            lcout => \FSM_TEST_inst_slow.counter_statZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10857\,
            ce => 'H',
            sr => \N__10638\
        );

    \FSM_TEST_inst_slow.counter_stat_4_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100011001001100"
        )
    port map (
            in0 => \N__9289\,
            in1 => \N__6029\,
            in2 => \N__9259\,
            in3 => \N__6035\,
            lcout => \FSM_TEST_inst_slow.counter_statZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10857\,
            ce => 'H',
            sr => \N__10638\
        );

    \FSM_TEST_inst_RAPIDA.current_state_RNO_0_0_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6008\,
            in1 => \N__5985\,
            in2 => \N__8463\,
            in3 => \N__5963\,
            lcout => \FSM_TEST_inst_RAPIDA.G_24_0_a4_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_RNI2J9G_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8455\,
            in2 => \_gnd_net_\,
            in3 => \N__11193\,
            lcout => \FSM_TEST_inst_RAPIDA.N_126_1_i\,
            ltout => \FSM_TEST_inst_RAPIDA.N_126_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_idle_1_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011011001100"
        )
    port map (
            in0 => \N__5942\,
            in1 => \N__6459\,
            in2 => \N__5933\,
            in3 => \N__6520\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10864\,
            ce => 'H',
            sr => \N__10635\
        );

    \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_RNI2J9G_0_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8454\,
            in2 => \_gnd_net_\,
            in3 => \N__11194\,
            lcout => \FSM_TEST_inst_RAPIDA.current_state_d_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.flag_output_1_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__11195\,
            in1 => \N__8462\,
            in2 => \N__11657\,
            in3 => \N__8061\,
            lcout => flag_signal,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10864\,
            ce => 'H',
            sr => \N__10635\
        );

    \FSM_TEST_inst_slow.flag_input_reg_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8062\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \FSM_TEST_inst_slow.flag_input_regZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10864\,
            ce => 'H',
            sr => \N__10635\
        );

    \FSM_TEST_inst_slow.current_state_RNO_4_0_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__7620\,
            in1 => \N__6210\,
            in2 => \N__6194\,
            in3 => \N__8768\,
            lcout => OPEN,
            ltout => \FSM_TEST_inst_slow.current_state_RNO_4Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.current_state_RNO_0_0_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__6184\,
            in1 => \N__6158\,
            in2 => \N__6152\,
            in3 => \N__6149\,
            lcout => \FSM_TEST_inst_slow.N_134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.current_state_RNO_3_0_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6335\,
            in1 => \N__11651\,
            in2 => \N__8468\,
            in3 => \N__6404\,
            lcout => \FSM_TEST_inst_RAPIDA.N_18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_0_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8467\,
            in2 => \_gnd_net_\,
            in3 => \N__11262\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10870\,
            ce => \N__12152\,
            sr => \N__10630\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_1_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11259\,
            in1 => \N__10330\,
            in2 => \_gnd_net_\,
            in3 => \N__6143\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10870\,
            ce => \N__12152\,
            sr => \N__10630\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_2_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11861\,
            in1 => \N__6137\,
            in2 => \_gnd_net_\,
            in3 => \N__11263\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10870\,
            ce => \N__12152\,
            sr => \N__10630\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_3_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11260\,
            in1 => \N__10331\,
            in2 => \_gnd_net_\,
            in3 => \N__6131\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10870\,
            ce => \N__12152\,
            sr => \N__10630\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_4_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10332\,
            in1 => \N__6365\,
            in2 => \_gnd_net_\,
            in3 => \N__11264\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10870\,
            ce => \N__12152\,
            sr => \N__10630\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_5_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11261\,
            in1 => \N__10333\,
            in2 => \_gnd_net_\,
            in3 => \N__6359\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10870\,
            ce => \N__12152\,
            sr => \N__10630\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_6_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11862\,
            in1 => \N__6353\,
            in2 => \_gnd_net_\,
            in3 => \N__11265\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10870\,
            ce => \N__12152\,
            sr => \N__10630\
        );

    \FSM_TEST_inst_RAPIDA.counter_idle_4_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001101000101010"
        )
    port map (
            in0 => \N__6316\,
            in1 => \N__6488\,
            in2 => \N__6530\,
            in3 => \N__6347\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10877\,
            ce => 'H',
            sr => \N__10625\
        );

    \FSM_TEST_inst_RAPIDA.current_state_RNO_6_0_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6294\,
            in1 => \N__6315\,
            in2 => \N__6277\,
            in3 => \N__6341\,
            lcout => \FSM_TEST_inst_RAPIDA.G_24_0_a4_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_idle_2_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001111100100000"
        )
    port map (
            in0 => \N__6329\,
            in1 => \N__6487\,
            in2 => \N__6529\,
            in3 => \N__6438\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10877\,
            ce => 'H',
            sr => \N__10625\
        );

    \FSM_TEST_inst_RAPIDA.counter_idle_3_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011010001110000"
        )
    port map (
            in0 => \N__6485\,
            in1 => \N__6521\,
            in2 => \N__6299\,
            in3 => \N__6323\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10877\,
            ce => 'H',
            sr => \N__10625\
        );

    \FSM_TEST_inst_RAPIDA.counter_idle_RNI23T81_5_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6314\,
            in1 => \N__6293\,
            in2 => \N__6278\,
            in3 => \N__6434\,
            lcout => OPEN,
            ltout => \FSM_TEST_inst_RAPIDA.counter_idlelde_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2_1_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__11271\,
            in1 => \N__9420\,
            in2 => \N__6533\,
            in3 => \N__11650\,
            lcout => \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1\,
            ltout => \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_idle_0_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101001101010"
        )
    port map (
            in0 => \N__6419\,
            in1 => \N__6609\,
            in2 => \N__6491\,
            in3 => \N__6486\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10877\,
            ce => 'H',
            sr => \N__10625\
        );

    \FSM_TEST_inst_RAPIDA.current_state_RNO_7_0_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__11270\,
            in1 => \N__6461\,
            in2 => \N__6440\,
            in3 => \N__6418\,
            lcout => \FSM_TEST_inst_RAPIDA.G_24_0_a4_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_7_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11282\,
            in1 => \N__10340\,
            in2 => \_gnd_net_\,
            in3 => \N__6398\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10883\,
            ce => \N__12151\,
            sr => \N__10620\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_19_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10334\,
            in1 => \N__7112\,
            in2 => \_gnd_net_\,
            in3 => \N__11283\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10883\,
            ce => \N__12151\,
            sr => \N__10620\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_20_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11279\,
            in1 => \N__10335\,
            in2 => \_gnd_net_\,
            in3 => \N__6389\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10883\,
            ce => \N__12151\,
            sr => \N__10620\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_21_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10336\,
            in1 => \N__6383\,
            in2 => \_gnd_net_\,
            in3 => \N__11284\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10883\,
            ce => \N__12151\,
            sr => \N__10620\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_22_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11280\,
            in1 => \N__10337\,
            in2 => \_gnd_net_\,
            in3 => \N__6377\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10883\,
            ce => \N__12151\,
            sr => \N__10620\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_23_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11281\,
            in1 => \N__10338\,
            in2 => \_gnd_net_\,
            in3 => \N__6371\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10883\,
            ce => \N__12151\,
            sr => \N__10620\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_24_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10339\,
            in1 => \N__6623\,
            in2 => \_gnd_net_\,
            in3 => \N__11285\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10883\,
            ce => \N__12151\,
            sr => \N__10620\
        );

    \CONSTANT_ONE_LUT4_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_86_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__6563\,
            in1 => \N__7811\,
            in2 => \_gnd_net_\,
            in3 => \N__9044\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10819\,
            ce => \N__7334\,
            sr => \N__10667\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_84_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__6551\,
            in1 => \N__7807\,
            in2 => \_gnd_net_\,
            in3 => \N__9042\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10820\,
            ce => \N__7333\,
            sr => \N__10663\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_85_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__9043\,
            in1 => \_gnd_net_\,
            in2 => \N__7915\,
            in3 => \N__6569\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10820\,
            ce => \N__7333\,
            sr => \N__10663\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_83_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__8979\,
            in1 => \_gnd_net_\,
            in2 => \N__7914\,
            in3 => \N__6557\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10822\,
            ce => \N__7332\,
            sr => \N__10658\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_12_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__6662\,
            in1 => \N__7800\,
            in2 => \_gnd_net_\,
            in3 => \N__8977\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10822\,
            ce => \N__7332\,
            sr => \N__10658\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_53_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__8978\,
            in1 => \_gnd_net_\,
            in2 => \N__7913\,
            in3 => \N__6539\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10822\,
            ce => \N__7332\,
            sr => \N__10658\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_7_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__6770\,
            in1 => \N__7781\,
            in2 => \_gnd_net_\,
            in3 => \N__8968\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10824\,
            ce => \N__7329\,
            sr => \N__10653\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_52_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110100101"
        )
    port map (
            in0 => \N__8966\,
            in1 => \_gnd_net_\,
            in2 => \N__7904\,
            in3 => \N__6635\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10824\,
            ce => \N__7329\,
            sr => \N__10653\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_10_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__6680\,
            in1 => \N__7773\,
            in2 => \_gnd_net_\,
            in3 => \N__8964\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10824\,
            ce => \N__7329\,
            sr => \N__10653\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_8_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110100101"
        )
    port map (
            in0 => \N__8969\,
            in1 => \_gnd_net_\,
            in2 => \N__7906\,
            in3 => \N__6692\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10824\,
            ce => \N__7329\,
            sr => \N__10653\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_9_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__6686\,
            in1 => \N__7785\,
            in2 => \_gnd_net_\,
            in3 => \N__8970\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10824\,
            ce => \N__7329\,
            sr => \N__10653\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_54_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__8967\,
            in1 => \_gnd_net_\,
            in2 => \N__7905\,
            in3 => \N__6674\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10824\,
            ce => \N__7329\,
            sr => \N__10653\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_11_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__6668\,
            in1 => \N__7774\,
            in2 => \_gnd_net_\,
            in3 => \N__8965\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10824\,
            ce => \N__7329\,
            sr => \N__10653\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_55_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__6656\,
            in1 => \N__7753\,
            in2 => \_gnd_net_\,
            in3 => \N__8960\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10828\,
            ce => \N__7326\,
            sr => \N__10649\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_56_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__8961\,
            in1 => \_gnd_net_\,
            in2 => \N__7899\,
            in3 => \N__6650\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10828\,
            ce => \N__7326\,
            sr => \N__10649\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_51_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__6644\,
            in1 => \N__7752\,
            in2 => \_gnd_net_\,
            in3 => \N__8959\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10828\,
            ce => \N__7326\,
            sr => \N__10649\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_6_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110100101"
        )
    port map (
            in0 => \N__8963\,
            in1 => \_gnd_net_\,
            in2 => \N__7900\,
            in3 => \N__6629\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10828\,
            ce => \N__7326\,
            sr => \N__10649\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_57_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__6764\,
            in1 => \N__7757\,
            in2 => \_gnd_net_\,
            in3 => \N__8962\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10828\,
            ce => \N__7326\,
            sr => \N__10649\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_69_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__6752\,
            in1 => \N__7536\,
            in2 => \_gnd_net_\,
            in3 => \N__8712\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10834\,
            ce => \N__7322\,
            sr => \N__10644\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_68_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__6746\,
            in1 => \N__7535\,
            in2 => \_gnd_net_\,
            in3 => \N__8711\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10834\,
            ce => \N__7322\,
            sr => \N__10644\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_67_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__7130\,
            in1 => \N__7534\,
            in2 => \_gnd_net_\,
            in3 => \N__8710\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10834\,
            ce => \N__7322\,
            sr => \N__10644\
        );

    \FSM_TEST_inst_slow.current_state_RNO_0_1_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8651\,
            in1 => \N__6943\,
            in2 => \N__6916\,
            in3 => \N__6891\,
            lcout => \FSM_TEST_inst_slow.current_state_cnv_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.current_state_RNIV6JP_1_1_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7457\,
            in2 => \_gnd_net_\,
            in3 => \N__8650\,
            lcout => \FSM_TEST_inst_slow.N_108_li\,
            ltout => \FSM_TEST_inst_slow.N_108_li_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.current_state_RNIR2L81_0_1_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6740\,
            in3 => \N__7208\,
            lcout => \FSM_TEST_inst_slow.current_state_RNIR2L81_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.current_state_1_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__7210\,
            in1 => \N__6725\,
            in2 => \_gnd_net_\,
            in3 => \N__7459\,
            lcout => \FSM_TEST_inst_slow.current_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10843\,
            ce => 'H',
            sr => \N__10639\
        );

    \FSM_TEST_inst_slow.counter_din_2_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110000010101010"
        )
    port map (
            in0 => \N__6912\,
            in1 => \N__6893\,
            in2 => \N__6716\,
            in3 => \N__7211\,
            lcout => \FSM_TEST_inst_slow.counter_dinZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10843\,
            ce => 'H',
            sr => \N__10639\
        );

    \FSM_TEST_inst_slow.current_state_RNO_8_0_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6944\,
            in1 => \N__6908\,
            in2 => \_gnd_net_\,
            in3 => \N__7458\,
            lcout => OPEN,
            ltout => \FSM_TEST_inst_slow.current_state_RNO_8Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.current_state_RNO_2_0_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101011111111"
        )
    port map (
            in0 => \N__8652\,
            in1 => \N__6892\,
            in2 => \N__6875\,
            in3 => \N__7209\,
            lcout => OPEN,
            ltout => \FSM_TEST_inst_slow.current_state_RNO_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.current_state_0_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110100001101"
        )
    port map (
            in0 => \N__6872\,
            in1 => \N__6866\,
            in2 => \N__6857\,
            in3 => \N__8653\,
            lcout => \FSM_TEST_inst_slow.current_stateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10843\,
            ce => 'H',
            sr => \N__10639\
        );

    \config_register_latched_dec_inst.DYNCNF_1_RNI9I121_8_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__9536\,
            in1 => \N__6832\,
            in2 => \N__12083\,
            in3 => \N__10098\,
            lcout => s12_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst.DYNCNF_1_8_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__9535\,
            in1 => \N__12063\,
            in2 => \N__6833\,
            in3 => \N__10085\,
            lcout => \config_register_latched_dec_inst.DYNCNF_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10851\,
            ce => \N__8078\,
            sr => \N__10636\
        );

    \config_register_latched_dec_inst.DYNCNF_1_9_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__10086\,
            in1 => \N__9505\,
            in2 => \N__12082\,
            in3 => \N__6820\,
            lcout => \config_register_latched_dec_inst.DYNCNF_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10851\,
            ce => \N__8078\,
            sr => \N__10636\
        );

    \config_register_latched_dec_inst.DYNCNF_1_RNIBK121_9_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__6821\,
            in1 => \N__12070\,
            in2 => \N__9509\,
            in3 => \N__10088\,
            lcout => s13_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst.DYNCNF_1_0_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__10087\,
            in1 => \N__8131\,
            in2 => \N__12081\,
            in3 => \N__6799\,
            lcout => \config_register_latched_dec_inst.DYNCNF_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10851\,
            ce => \N__8078\,
            sr => \N__10636\
        );

    \config_register_latched_dec_inst.DYNCNF_1_RNIP1121_0_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010100000"
        )
    port map (
            in0 => \N__6800\,
            in1 => \N__12071\,
            in2 => \N__10105\,
            in3 => \N__8132\,
            lcout => \config_register_latched_dec_inst.DYNCNF_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst.DYNCNF_1_10_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__8179\,
            in1 => \N__12062\,
            in2 => \N__8002\,
            in3 => \N__10084\,
            lcout => \config_register_latched_dec_inst.DYNCNF_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10851\,
            ce => \N__8078\,
            sr => \N__10636\
        );

    \FSM_TEST_inst_RAPIDA.counter_din_RNO_0_2_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__9932\,
            in1 => \N__9879\,
            in2 => \N__9977\,
            in3 => \N__11908\,
            lcout => OPEN,
            ltout => \FSM_TEST_inst_RAPIDA.counter_din_3_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_din_2_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__9971\,
            in1 => \N__8191\,
            in2 => \N__7040\,
            in3 => \N__11616\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10858\,
            ce => 'H',
            sr => \N__10631\
        );

    \FSM_TEST_inst_RAPIDA.current_state_RNO_5_0_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__9931\,
            in1 => \N__9970\,
            in2 => \N__9909\,
            in3 => \N__9878\,
            lcout => OPEN,
            ltout => \FSM_TEST_inst_RAPIDA.G_24_0_o4_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.current_state_RNO_2_0_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__8456\,
            in1 => \N__11613\,
            in2 => \N__7037\,
            in3 => \N__11220\,
            lcout => \FSM_TEST_inst_RAPIDA.N_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.current_state_RNO_1_0_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__11614\,
            in1 => \N__7034\,
            in2 => \N__7025\,
            in3 => \N__6992\,
            lcout => OPEN,
            ltout => \FSM_TEST_inst_RAPIDA.G_24_0_a4_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.current_state_0_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__6965\,
            in1 => \N__6959\,
            in2 => \N__6953\,
            in3 => \N__6950\,
            lcout => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10858\,
            ce => 'H',
            sr => \N__10631\
        );

    \FSM_TEST_inst_RAPIDA.counter_din_1_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100001010000"
        )
    port map (
            in0 => \N__11615\,
            in1 => \N__9880\,
            in2 => \N__9940\,
            in3 => \N__11909\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_dinZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10858\,
            ce => 'H',
            sr => \N__10631\
        );

    \FSM_TEST_inst_RAPIDA.counter_din_3_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100011110000"
        )
    port map (
            in0 => \N__11910\,
            in1 => \N__8192\,
            in2 => \N__9910\,
            in3 => \N__11617\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10858\,
            ce => 'H',
            sr => \N__10631\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_15_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11254\,
            in2 => \N__10341\,
            in3 => \N__7118\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10865\,
            ce => \N__8233\,
            sr => \N__10626\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_0_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__11258\,
            in1 => \N__9413\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10865\,
            ce => \N__8233\,
            sr => \N__10626\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_5_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11256\,
            in2 => \N__10342\,
            in3 => \N__7064\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10865\,
            ce => \N__8233\,
            sr => \N__10626\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_1_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__7076\,
            in1 => \N__9414\,
            in2 => \_gnd_net_\,
            in3 => \N__11266\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10865\,
            ce => \N__8233\,
            sr => \N__10626\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_2_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11255\,
            in2 => \N__9424\,
            in3 => \N__7070\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10865\,
            ce => \N__8233\,
            sr => \N__10626\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_4_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__7046\,
            in1 => \N__9419\,
            in2 => \_gnd_net_\,
            in3 => \N__11268\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10865\,
            ce => \N__8233\,
            sr => \N__10626\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_6_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11257\,
            in2 => \N__10343\,
            in3 => \N__7058\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10865\,
            ce => \N__8233\,
            sr => \N__10626\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_3_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__7052\,
            in1 => \N__9418\,
            in2 => \_gnd_net_\,
            in3 => \N__11267\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10865\,
            ce => \N__8233\,
            sr => \N__10626\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_13_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10324\,
            in1 => \N__8243\,
            in2 => \_gnd_net_\,
            in3 => \N__11286\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10871\,
            ce => \N__8237\,
            sr => \N__10621\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_14_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10325\,
            in1 => \N__7124\,
            in2 => \_gnd_net_\,
            in3 => \N__11287\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10871\,
            ce => \N__8237\,
            sr => \N__10621\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_18_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10326\,
            in1 => \N__9755\,
            in2 => \_gnd_net_\,
            in3 => \N__11275\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10878\,
            ce => \N__12149\,
            sr => \N__10615\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_79_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11045\,
            in1 => \N__7100\,
            in2 => \_gnd_net_\,
            in3 => \N__11278\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10878\,
            ce => \N__12149\,
            sr => \N__10615\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_27_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11273\,
            in1 => \N__10328\,
            in2 => \_gnd_net_\,
            in3 => \N__7082\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10878\,
            ce => \N__12149\,
            sr => \N__10615\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_25_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__7106\,
            in1 => \N__10329\,
            in2 => \_gnd_net_\,
            in3 => \N__11276\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10878\,
            ce => \N__12149\,
            sr => \N__10615\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_78_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11274\,
            in1 => \N__11044\,
            in2 => \_gnd_net_\,
            in3 => \N__7094\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10878\,
            ce => \N__12149\,
            sr => \N__10615\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_77_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11864\,
            in1 => \N__8408\,
            in2 => \_gnd_net_\,
            in3 => \N__11277\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10878\,
            ce => \N__12149\,
            sr => \N__10615\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_26_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11272\,
            in1 => \N__10327\,
            in2 => \_gnd_net_\,
            in3 => \N__7088\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10878\,
            ce => \N__12149\,
            sr => \N__10615\
        );

    \FSM_TEST_inst_RAPIDA.CLK_uC_4_0_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7184\,
            lcout => \FSM_TEST_inst_RAPIDA.CLK_uC_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10884\,
            ce => 'H',
            sr => \N__10611\
        );

    \FSM_TEST_inst_RAPIDA.CLK_uC_6_0_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7172\,
            lcout => \FSM_TEST_inst_RAPIDA.CLK_uC_6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10884\,
            ce => 'H',
            sr => \N__10611\
        );

    \FSM_TEST_inst_RAPIDA.CLK_uC_3_0_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8396\,
            lcout => \FSM_TEST_inst_RAPIDA.CLK_uC_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10884\,
            ce => 'H',
            sr => \N__10611\
        );

    \FSM_TEST_inst_RAPIDA.CLK_uC_5_0_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7178\,
            lcout => \FSM_TEST_inst_RAPIDA.CLK_uC_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10884\,
            ce => 'H',
            sr => \N__10611\
        );

    \FSM_TEST_inst_RAPIDA.CLK_uC_6b_0_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7166\,
            lcout => \FSM_TEST_inst_RAPIDA.CLK_uC_6bZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10884\,
            ce => 'H',
            sr => \N__10611\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_61_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__8941\,
            in1 => \N__7154\,
            in2 => \_gnd_net_\,
            in3 => \N__7799\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10825\,
            ce => \N__7330\,
            sr => \N__10645\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_58_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__7796\,
            in1 => \N__7160\,
            in2 => \_gnd_net_\,
            in3 => \N__8938\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10825\,
            ce => \N__7330\,
            sr => \N__10645\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_60_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__8940\,
            in1 => \N__7142\,
            in2 => \_gnd_net_\,
            in3 => \N__7798\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10825\,
            ce => \N__7330\,
            sr => \N__10645\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_59_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__8939\,
            in1 => \N__7148\,
            in2 => \_gnd_net_\,
            in3 => \N__7797\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10825\,
            ce => \N__7330\,
            sr => \N__10645\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_62_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__7136\,
            in1 => \N__7568\,
            in2 => \_gnd_net_\,
            in3 => \N__8720\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10829\,
            ce => \N__7327\,
            sr => \N__10640\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_66_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__8724\,
            in1 => \N__7952\,
            in2 => \_gnd_net_\,
            in3 => \N__7572\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10829\,
            ce => \N__7327\,
            sr => \N__10640\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_64_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__7340\,
            in1 => \N__7569\,
            in2 => \_gnd_net_\,
            in3 => \N__8722\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10829\,
            ce => \N__7327\,
            sr => \N__10640\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_65_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__8723\,
            in1 => \N__7958\,
            in2 => \_gnd_net_\,
            in3 => \N__7571\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10829\,
            ce => \N__7327\,
            sr => \N__10640\
        );

    \FSM_TEST_inst_slow.bit_sequence_stat_63_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__8721\,
            in1 => \N__7946\,
            in2 => \_gnd_net_\,
            in3 => \N__7570\,
            lcout => \FSM_TEST_inst_slow.bit_sequence_statZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10829\,
            ce => \N__7327\,
            sr => \N__10640\
        );

    \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5D1_0_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__11598\,
            in1 => \N__8496\,
            in2 => \N__9085\,
            in3 => \N__11269\,
            lcout => \N_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divisor_inst_2.counter_RNIFD27_2_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__9163\,
            in1 => \_gnd_net_\,
            in2 => \N__9110\,
            in3 => \N__9130\,
            lcout => \counter_RNIFD27_2\,
            ltout => \counter_RNIFD27_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_slow.SEL_0_RNI25J31_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__8534\,
            in1 => \N__8513\,
            in2 => \N__7253\,
            in3 => \N__8709\,
            lcout => \N_3_0\,
            ltout => \N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst.STATCNF_1_RNO_0_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8351\,
            in2 => \N__7250\,
            in3 => \N__7247\,
            lcout => \config_register_latched_dec_inst.N_378_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divisor_inst_2.counter_RNISR1F_2_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__9162\,
            in1 => \N__9129\,
            in2 => \N__9109\,
            in3 => \N__8533\,
            lcout => \counter_RNISR1F_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divisor_inst_2.clk_out_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__8535\,
            in1 => \N__9164\,
            in2 => \N__9139\,
            in3 => \N__9107\,
            lcout => clk_continuous_slow,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10835\,
            ce => 'H',
            sr => \N__10637\
        );

    \FSM_TEST_inst_RAPIDA.MOSI_er_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000010001000"
        )
    port map (
            in0 => \N__11149\,
            in1 => \N__8099\,
            in2 => \N__9671\,
            in3 => \N__8433\,
            lcout => mosi_fast,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10844\,
            ce => \N__11642\,
            sr => \N__10632\
        );

    \divisor_inst.clk_out_RNI3LEM_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__11992\,
            in1 => \N__11930\,
            in2 => \_gnd_net_\,
            in3 => \N__11960\,
            lcout => \clk_out_RNI3LEM\,
            ltout => \clk_out_RNI3LEM_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.flag_output_1_RNIVLAE1_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__11148\,
            in1 => \N__8068\,
            in2 => \N__8087\,
            in3 => \N__8432\,
            lcout => \N_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIHTFF_1_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8486\,
            in2 => \_gnd_net_\,
            in3 => \N__11147\,
            lcout => \FSM_TEST_inst_RAPIDA.N_100_li\,
            ltout => \FSM_TEST_inst_RAPIDA.N_100_li_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5D1_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9081\,
            in2 => \N__8084\,
            in3 => \N__11599\,
            lcout => \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5DZ0Z1\,
            ltout => \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5DZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.SEL_0_RNI8H3V3_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__8365\,
            in1 => \_gnd_net_\,
            in2 => \N__8081\,
            in3 => \N__8350\,
            lcout => \N_378_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mosi_output_obuf_RNO_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8069\,
            in1 => \N__8045\,
            in2 => \_gnd_net_\,
            in3 => \N__8039\,
            lcout => mosi_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst.DYNCNF_1_RNIR83V_10_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__10082\,
            in1 => \N__12095\,
            in2 => \N__8180\,
            in3 => \N__8003\,
            lcout => s14_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst.STATCNF_1_0_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__10081\,
            in1 => \N__12096\,
            in2 => \N__10153\,
            in3 => \N__10123\,
            lcout => \config_register_latched_dec_inst.STATCNF_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10852\,
            ce => \N__7967\,
            sr => \N__10627\
        );

    \flag_output_0_ret_RNI1E8N2_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__9343\,
            in1 => \N__8290\,
            in2 => \N__8326\,
            in3 => \N__8352\,
            lcout => \flag_output_0_ret_RNI1E8NZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_din_RNI9NO1_1_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9973\,
            in1 => \N__9936\,
            in2 => \_gnd_net_\,
            in3 => \N__9873\,
            lcout => \FSM_TEST_inst_RAPIDA.N_101_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.current_state_fast_RNI78E11_1_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__9387\,
            in1 => \N__11618\,
            in2 => \_gnd_net_\,
            in3 => \N__11219\,
            lcout => \FSM_TEST_inst_RAPIDA.current_state_fast_RNI78E11Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst.DYNSR_10_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10083\,
            in1 => \N__8175\,
            in2 => \_gnd_net_\,
            in3 => \N__9499\,
            lcout => \config_register_latched_dec_inst.DYNSRZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10859\,
            ce => \N__9478\,
            sr => \N__10622\
        );

    \config_register_latched_dec_inst.STATSR_0_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10079\,
            in1 => \N__8156\,
            in2 => \_gnd_net_\,
            in3 => \N__10149\,
            lcout => \config_register_latched_dec_inst.STATSRZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10859\,
            ce => \N__9478\,
            sr => \N__10622\
        );

    \config_register_latched_dec_inst.DYNSR_1_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8123\,
            in1 => \N__10080\,
            in2 => \_gnd_net_\,
            in3 => \N__9314\,
            lcout => \config_register_latched_dec_inst.DYNSRZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10859\,
            ce => \N__9478\,
            sr => \N__10622\
        );

    \config_register_latched_dec_inst.DYNSR_0_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10078\,
            in1 => \N__8155\,
            in2 => \_gnd_net_\,
            in3 => \N__8124\,
            lcout => \config_register_latched_dec_inst.DYNSRZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10859\,
            ce => \N__9478\,
            sr => \N__10622\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_10_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11481\,
            in1 => \N__8255\,
            in2 => \_gnd_net_\,
            in3 => \N__10245\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10866\,
            ce => \N__8232\,
            sr => \N__10616\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_11_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11477\,
            in2 => \N__10311\,
            in3 => \N__8105\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10866\,
            ce => \N__8232\,
            sr => \N__10616\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_8_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11480\,
            in2 => \N__10314\,
            in3 => \N__8267\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10866\,
            ce => \N__8232\,
            sr => \N__10616\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_7_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11479\,
            in2 => \N__10313\,
            in3 => \N__8273\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10866\,
            ce => \N__8232\,
            sr => \N__10616\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_9_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11482\,
            in1 => \N__8261\,
            in2 => \_gnd_net_\,
            in3 => \N__10258\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10866\,
            ce => \N__8232\,
            sr => \N__10616\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_din_12_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11478\,
            in2 => \N__10312\,
            in3 => \N__8249\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10866\,
            ce => \N__8232\,
            sr => \N__10616\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_59_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11041\,
            in1 => \N__9608\,
            in2 => \_gnd_net_\,
            in3 => \N__11488\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10872\,
            ce => \N__12146\,
            sr => \N__10612\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_54_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11483\,
            in1 => \N__11040\,
            in2 => \_gnd_net_\,
            in3 => \N__9443\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10872\,
            ce => \N__12146\,
            sr => \N__10612\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_29_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10259\,
            in1 => \N__8204\,
            in2 => \_gnd_net_\,
            in3 => \N__11487\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10872\,
            ce => \N__12146\,
            sr => \N__10612\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_28_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11039\,
            in1 => \N__8210\,
            in2 => \_gnd_net_\,
            in3 => \N__11486\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10872\,
            ce => \N__12146\,
            sr => \N__10612\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_60_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11485\,
            in1 => \N__11042\,
            in2 => \_gnd_net_\,
            in3 => \N__8198\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10872\,
            ce => \N__12146\,
            sr => \N__10612\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_76_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11043\,
            in1 => \N__9620\,
            in2 => \_gnd_net_\,
            in3 => \N__11489\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10872\,
            ce => \N__12146\,
            sr => \N__10612\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_55_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11484\,
            in1 => \N__11863\,
            in2 => \_gnd_net_\,
            in3 => \N__8402\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10872\,
            ce => \N__12146\,
            sr => \N__10612\
        );

    \FSM_TEST_inst_RAPIDA.CLK_uC_2_0_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8383\,
            lcout => \FSM_TEST_inst_RAPIDA.CLK_uC_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10879\,
            ce => 'H',
            sr => \N__10608\
        );

    \FSM_TEST_inst_RAPIDA.CLK_uC_6c_0_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8390\,
            lcout => \CLK_uC_6c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10879\,
            ce => 'H',
            sr => \N__10608\
        );

    \FSM_TEST_inst_RAPIDA.CLK_uC_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011010010000"
        )
    port map (
            in0 => \N__11466\,
            in1 => \N__9425\,
            in2 => \N__8384\,
            in3 => \N__11972\,
            lcout => \FSM_TEST_inst_RAPIDA.CLK_uCZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10879\,
            ce => 'H',
            sr => \N__10608\
        );

    \flag_output_ret_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8372\,
            in1 => \N__8366\,
            in2 => \_gnd_net_\,
            in3 => \N__8353\,
            lcout => sel_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10830\,
            ce => 'H',
            sr => \N__10633\
        );

    \flag_output_0_ret_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8354\,
            in1 => \N__9347\,
            in2 => \_gnd_net_\,
            in3 => \N__8327\,
            lcout => clk_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10830\,
            ce => 'H',
            sr => \N__10633\
        );

    \divisor_inst_2.counter_1_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9134\,
            in2 => \_gnd_net_\,
            in3 => \N__9160\,
            lcout => \divisor_inst_2.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10830\,
            ce => 'H',
            sr => \N__10633\
        );

    \divisor_inst_2.counter_0_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9135\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \divisor_inst_2.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10830\,
            ce => 'H',
            sr => \N__10633\
        );

    \FSM_TEST_inst_slow.counter_stat_5_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100011001001100"
        )
    port map (
            in0 => \N__9292\,
            in1 => \N__9182\,
            in2 => \N__9260\,
            in3 => \N__9206\,
            lcout => \FSM_TEST_inst_slow.counter_statZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10830\,
            ce => 'H',
            sr => \N__10633\
        );

    \divisor_inst_2.counter_2_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110001101100"
        )
    port map (
            in0 => \N__9161\,
            in1 => \N__9108\,
            in2 => \N__9140\,
            in3 => \_gnd_net_\,
            lcout => \divisor_inst_2.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10830\,
            ce => 'H',
            sr => \N__10633\
        );

    \FSM_TEST_inst_RAPIDA.SEL_0_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__8497\,
            in1 => \N__11619\,
            in2 => \N__9086\,
            in3 => \N__11534\,
            lcout => \FSM_TEST_inst_RAPIDA.aux_selection_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10830\,
            ce => 'H',
            sr => \N__10633\
        );

    \FSM_TEST_inst_slow.SEL_0_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__8512\,
            in1 => \N__9012\,
            in2 => \N__8555\,
            in3 => \N__8536\,
            lcout => \FSM_TEST_inst_slow.aux_selection_slow_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10836\,
            ce => 'H',
            sr => \N__10628\
        );

    \divisor_inst.clk_out_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__11935\,
            in1 => \N__11998\,
            in2 => \_gnd_net_\,
            in3 => \N__11964\,
            lcout => clk_continuous_fast,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10836\,
            ce => 'H',
            sr => \N__10628\
        );

    \divisor_inst.counter_1_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11997\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11934\,
            lcout => divisor_inst_counter_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10836\,
            ce => 'H',
            sr => \N__10628\
        );

    \divisor_inst.counter_0_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11996\,
            lcout => divisor_inst_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10836\,
            ce => 'H',
            sr => \N__10628\
        );

    \FSM_TEST_inst_RAPIDA.current_state_fast_fast_1_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__11624\,
            in1 => \N__11369\,
            in2 => \N__8498\,
            in3 => \N__11689\,
            lcout => \FSM_TEST_inst_RAPIDA.current_state_fast_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10845\,
            ce => 'H',
            sr => \N__10623\
        );

    \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__11366\,
            in1 => \N__8450\,
            in2 => \N__11690\,
            in3 => \N__11623\,
            lcout => \FSM_TEST_inst_RAPIDA.current_state_fast_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10845\,
            ce => 'H',
            sr => \N__10623\
        );

    \FSM_TEST_inst_RAPIDA.current_state_fast_1_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__11622\,
            in1 => \N__11685\,
            in2 => \N__9411\,
            in3 => \N__11368\,
            lcout => \FSM_TEST_inst_RAPIDA.current_state_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10845\,
            ce => 'H',
            sr => \N__10623\
        );

    \FSM_TEST_inst_slow.CLK_uC_6l_0_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9356\,
            lcout => \CLK_uC_6l_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10845\,
            ce => 'H',
            sr => \N__10623\
        );

    \FSM_TEST_inst_RAPIDA.current_state_1_rep1_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__11621\,
            in1 => \N__11684\,
            in2 => \N__10243\,
            in3 => \N__11367\,
            lcout => \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10845\,
            ce => 'H',
            sr => \N__10623\
        );

    \FSM_TEST_inst_RAPIDA.counter_din_0_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011001000100"
        )
    port map (
            in0 => \N__11620\,
            in1 => \N__9877\,
            in2 => \_gnd_net_\,
            in3 => \N__11911\,
            lcout => \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10845\,
            ce => 'H',
            sr => \N__10623\
        );

    \config_register_latched_dec_inst.DYNSR_3_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9332\,
            in1 => \N__10073\,
            in2 => \_gnd_net_\,
            in3 => \N__9301\,
            lcout => \config_register_latched_dec_inst.DYNSRZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10853\,
            ce => \N__9479\,
            sr => \N__10617\
        );

    \config_register_latched_dec_inst.DYNSR_4_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9323\,
            in1 => \N__10069\,
            in2 => \_gnd_net_\,
            in3 => \N__9331\,
            lcout => \config_register_latched_dec_inst.DYNSRZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10853\,
            ce => \N__9479\,
            sr => \N__10617\
        );

    \config_register_latched_dec_inst.DYNSR_5_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10068\,
            in1 => \N__9554\,
            in2 => \_gnd_net_\,
            in3 => \N__9322\,
            lcout => \config_register_latched_dec_inst.DYNSRZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10853\,
            ce => \N__9479\,
            sr => \N__10617\
        );

    \config_register_latched_dec_inst.DYNSR_7_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10070\,
            in1 => \N__9563\,
            in2 => \_gnd_net_\,
            in3 => \N__9544\,
            lcout => \config_register_latched_dec_inst.DYNSRZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10853\,
            ce => \N__9479\,
            sr => \N__10617\
        );

    \config_register_latched_dec_inst.DYNSR_2_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10067\,
            in1 => \N__9302\,
            in2 => \_gnd_net_\,
            in3 => \N__9313\,
            lcout => \config_register_latched_dec_inst.DYNSRZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10853\,
            ce => \N__9479\,
            sr => \N__10617\
        );

    \config_register_latched_dec_inst.DYNSR_8_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10071\,
            in1 => \N__9527\,
            in2 => \_gnd_net_\,
            in3 => \N__9562\,
            lcout => \config_register_latched_dec_inst.DYNSRZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10853\,
            ce => \N__9479\,
            sr => \N__10617\
        );

    \config_register_latched_dec_inst.DYNSR_6_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9545\,
            in1 => \N__10074\,
            in2 => \_gnd_net_\,
            in3 => \N__9553\,
            lcout => \config_register_latched_dec_inst.DYNSRZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10853\,
            ce => \N__9479\,
            sr => \N__10617\
        );

    \config_register_latched_dec_inst.DYNSR_9_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10072\,
            in1 => \N__9498\,
            in2 => \_gnd_net_\,
            in3 => \N__9528\,
            lcout => \config_register_latched_dec_inst.DYNSRZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10853\,
            ce => \N__9479\,
            sr => \N__10617\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_31_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__9626\,
            in1 => \N__11847\,
            in2 => \_gnd_net_\,
            in3 => \N__11463\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10860\,
            ce => \N__12147\,
            sr => \N__10613\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_52_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11462\,
            in1 => \N__11030\,
            in2 => \_gnd_net_\,
            in3 => \N__9455\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10860\,
            ce => \N__12147\,
            sr => \N__10613\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_51_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11461\,
            in1 => \N__9431\,
            in2 => \_gnd_net_\,
            in3 => \N__11851\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10860\,
            ce => \N__12147\,
            sr => \N__10613\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_53_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11031\,
            in1 => \N__9449\,
            in2 => \_gnd_net_\,
            in3 => \N__11465\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10860\,
            ce => \N__12147\,
            sr => \N__10613\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_32_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11460\,
            in2 => \N__11870\,
            in3 => \N__9437\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10860\,
            ce => \N__12147\,
            sr => \N__10613\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_50_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11029\,
            in1 => \N__9809\,
            in2 => \_gnd_net_\,
            in3 => \N__11464\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10860\,
            ce => \N__12147\,
            sr => \N__10613\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_9_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11469\,
            in1 => \N__11869\,
            in2 => \_gnd_net_\,
            in3 => \N__9593\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10867\,
            ce => \N__12143\,
            sr => \N__10609\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_30_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11865\,
            in1 => \N__9632\,
            in2 => \_gnd_net_\,
            in3 => \N__11471\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10867\,
            ce => \N__12143\,
            sr => \N__10609\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_75_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11033\,
            in1 => \N__9785\,
            in2 => \_gnd_net_\,
            in3 => \N__11473\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10867\,
            ce => \N__12143\,
            sr => \N__10609\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_61_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11467\,
            in1 => \N__11867\,
            in2 => \_gnd_net_\,
            in3 => \N__9614\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10867\,
            ce => \N__12143\,
            sr => \N__10609\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_58_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11866\,
            in1 => \N__9581\,
            in2 => \_gnd_net_\,
            in3 => \N__11472\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10867\,
            ce => \N__12143\,
            sr => \N__10609\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_8_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11468\,
            in1 => \N__11868\,
            in2 => \_gnd_net_\,
            in3 => \N__9602\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10867\,
            ce => \N__12143\,
            sr => \N__10609\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_10_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10244\,
            in1 => \N__9587\,
            in2 => \_gnd_net_\,
            in3 => \N__11470\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10867\,
            ce => \N__12143\,
            sr => \N__10609\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_57_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11474\,
            in1 => \N__11872\,
            in2 => \_gnd_net_\,
            in3 => \N__9683\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10873\,
            ce => \N__12140\,
            sr => \N__10605\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_80_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11475\,
            in1 => \N__11873\,
            in2 => \_gnd_net_\,
            in3 => \N__9575\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10873\,
            ce => \N__12140\,
            sr => \N__10605\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_56_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11871\,
            in1 => \N__9689\,
            in2 => \_gnd_net_\,
            in3 => \N__11476\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10873\,
            ce => \N__12140\,
            sr => \N__10605\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_83_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10968\,
            in1 => \N__9638\,
            in2 => \_gnd_net_\,
            in3 => \N__11456\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10837\,
            ce => \N__12150\,
            sr => \N__10618\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_84_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11454\,
            in1 => \N__10969\,
            in2 => \_gnd_net_\,
            in3 => \N__9677\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10837\,
            ce => \N__12150\,
            sr => \N__10618\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_87_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10972\,
            in1 => \N__9644\,
            in2 => \_gnd_net_\,
            in3 => \N__11458\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10837\,
            ce => \N__12150\,
            sr => \N__10618\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_85_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10970\,
            in1 => \N__9656\,
            in2 => \_gnd_net_\,
            in3 => \N__11457\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10837\,
            ce => \N__12150\,
            sr => \N__10618\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_86_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11455\,
            in1 => \N__10971\,
            in2 => \_gnd_net_\,
            in3 => \N__9650\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10837\,
            ce => \N__12150\,
            sr => \N__10618\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_46_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11496\,
            in1 => \N__11023\,
            in2 => \_gnd_net_\,
            in3 => \N__9833\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10846\,
            ce => \N__12148\,
            sr => \N__10614\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_35_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11810\,
            in1 => \N__9797\,
            in2 => \_gnd_net_\,
            in3 => \N__11498\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10846\,
            ce => \N__12148\,
            sr => \N__10614\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_82_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11025\,
            in1 => \N__9725\,
            in2 => \_gnd_net_\,
            in3 => \N__11501\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10846\,
            ce => \N__12148\,
            sr => \N__10614\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_66_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11497\,
            in1 => \N__11812\,
            in2 => \_gnd_net_\,
            in3 => \N__9746\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10846\,
            ce => \N__12148\,
            sr => \N__10614\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_65_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11024\,
            in1 => \N__10406\,
            in2 => \_gnd_net_\,
            in3 => \N__11500\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10846\,
            ce => \N__12148\,
            sr => \N__10614\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_36_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11495\,
            in1 => \N__11022\,
            in2 => \_gnd_net_\,
            in3 => \N__9740\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10846\,
            ce => \N__12148\,
            sr => \N__10614\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_40_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11811\,
            in1 => \N__9713\,
            in2 => \_gnd_net_\,
            in3 => \N__11499\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10846\,
            ce => \N__12148\,
            sr => \N__10614\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_81_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11505\,
            in1 => \N__11028\,
            in2 => \_gnd_net_\,
            in3 => \N__9734\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10854\,
            ce => \N__12144\,
            sr => \N__10610\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_33_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11026\,
            in1 => \N__9719\,
            in2 => \_gnd_net_\,
            in3 => \N__11506\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10854\,
            ce => \N__12144\,
            sr => \N__10610\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_39_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11502\,
            in1 => \N__11832\,
            in2 => \_gnd_net_\,
            in3 => \N__9827\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10854\,
            ce => \N__12144\,
            sr => \N__10610\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_48_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11835\,
            in1 => \N__9701\,
            in2 => \_gnd_net_\,
            in3 => \N__11509\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10854\,
            ce => \N__12144\,
            sr => \N__10610\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_47_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11503\,
            in1 => \N__11834\,
            in2 => \_gnd_net_\,
            in3 => \N__9707\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10854\,
            ce => \N__12144\,
            sr => \N__10610\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_41_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11833\,
            in1 => \N__9695\,
            in2 => \_gnd_net_\,
            in3 => \N__11508\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10854\,
            ce => \N__12144\,
            sr => \N__10610\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_49_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11504\,
            in1 => \N__11027\,
            in2 => \_gnd_net_\,
            in3 => \N__9815\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10854\,
            ce => \N__12144\,
            sr => \N__10610\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_34_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11831\,
            in1 => \N__9803\,
            in2 => \_gnd_net_\,
            in3 => \N__11507\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10854\,
            ce => \N__12144\,
            sr => \N__10610\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_11_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11513\,
            in1 => \N__10306\,
            in2 => \_gnd_net_\,
            in3 => \N__9791\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10861\,
            ce => \N__12141\,
            sr => \N__10606\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_74_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__12158\,
            in1 => \N__11032\,
            in2 => \_gnd_net_\,
            in3 => \N__11520\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10861\,
            ce => \N__12141\,
            sr => \N__10606\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_16_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11515\,
            in1 => \N__11853\,
            in2 => \_gnd_net_\,
            in3 => \N__9767\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10861\,
            ce => \N__12141\,
            sr => \N__10606\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_13_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11852\,
            in1 => \N__10163\,
            in2 => \_gnd_net_\,
            in3 => \N__11518\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10861\,
            ce => \N__12141\,
            sr => \N__10606\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_14_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11514\,
            in1 => \N__10308\,
            in2 => \_gnd_net_\,
            in3 => \N__9779\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10861\,
            ce => \N__12141\,
            sr => \N__10606\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_15_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10309\,
            in1 => \N__9773\,
            in2 => \_gnd_net_\,
            in3 => \N__11519\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10861\,
            ce => \N__12141\,
            sr => \N__10606\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_17_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11516\,
            in1 => \N__10310\,
            in2 => \_gnd_net_\,
            in3 => \N__9761\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10861\,
            ce => \N__12141\,
            sr => \N__10606\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_12_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10307\,
            in1 => \N__10169\,
            in2 => \_gnd_net_\,
            in3 => \N__11517\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10861\,
            ce => \N__12141\,
            sr => \N__10606\
        );

    \config_register_latched_dec_inst.STATCNF_1_RNIRDN51_0_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__12097\,
            in1 => \N__10157\,
            in2 => \N__10130\,
            in3 => \N__10094\,
            lcout => \config_register_latched_dec_inst.STATCNF_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.counter_din_RNIEMB2_3_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9972\,
            in1 => \N__9941\,
            in2 => \N__9911\,
            in3 => \N__9881\,
            lcout => \FSM_TEST_inst_RAPIDA.N_123_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_68_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10944\,
            in1 => \N__9839\,
            in2 => \_gnd_net_\,
            in3 => \N__11512\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10831\,
            ce => \N__12145\,
            sr => \N__10607\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_67_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11510\,
            in1 => \N__10943\,
            in2 => \_gnd_net_\,
            in3 => \N__9845\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10831\,
            ce => \N__12145\,
            sr => \N__10607\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_45_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11723\,
            in1 => \N__10412\,
            in2 => \_gnd_net_\,
            in3 => \N__11511\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10831\,
            ce => \N__12145\,
            sr => \N__10607\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_38_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11521\,
            in1 => \N__11824\,
            in2 => \_gnd_net_\,
            in3 => \N__10424\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10840\,
            ce => \N__12142\,
            sr => \N__10604\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_43_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__11522\,
            in1 => \_gnd_net_\,
            in2 => \N__10364\,
            in3 => \N__11825\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10840\,
            ce => \N__12142\,
            sr => \N__10604\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_37_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10999\,
            in1 => \N__9821\,
            in2 => \_gnd_net_\,
            in3 => \N__11524\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10840\,
            ce => \N__12142\,
            sr => \N__10604\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_44_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11000\,
            in1 => \N__10418\,
            in2 => \_gnd_net_\,
            in3 => \N__11525\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10840\,
            ce => \N__12142\,
            sr => \N__10604\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_64_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11523\,
            in1 => \N__11826\,
            in2 => \_gnd_net_\,
            in3 => \N__10400\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10840\,
            ce => \N__12142\,
            sr => \N__10604\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_63_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11001\,
            in1 => \N__10385\,
            in2 => \_gnd_net_\,
            in3 => \N__11526\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10840\,
            ce => \N__12142\,
            sr => \N__10604\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_62_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11827\,
            in1 => \N__10394\,
            in2 => \_gnd_net_\,
            in3 => \N__11531\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10848\,
            ce => \N__12139\,
            sr => \N__10603\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_69_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__11527\,
            in1 => \N__11003\,
            in2 => \_gnd_net_\,
            in3 => \N__10379\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10848\,
            ce => \N__12139\,
            sr => \N__10603\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_42_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11002\,
            in1 => \N__10370\,
            in2 => \_gnd_net_\,
            in3 => \N__11530\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10848\,
            ce => \N__12139\,
            sr => \N__10603\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_70_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11528\,
            in1 => \N__11828\,
            in2 => \_gnd_net_\,
            in3 => \N__10355\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10848\,
            ce => \N__12139\,
            sr => \N__10603\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_71_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__11004\,
            in1 => \N__10349\,
            in2 => \_gnd_net_\,
            in3 => \N__11532\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10848\,
            ce => \N__12139\,
            sr => \N__10603\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_72_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11529\,
            in1 => \N__11829\,
            in2 => \_gnd_net_\,
            in3 => \N__12170\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10848\,
            ce => \N__12139\,
            sr => \N__10603\
        );

    \FSM_TEST_inst_RAPIDA.bit_sequence_stat_73_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11830\,
            in1 => \N__12164\,
            in2 => \_gnd_net_\,
            in3 => \N__11533\,
            lcout => \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10848\,
            ce => \N__12139\,
            sr => \N__10603\
        );

    \RST_N_ibuf_RNIBJGC_LC_16_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12034\,
            lcout => \RST_N_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIKIU51_1_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__11999\,
            in1 => \N__11968\,
            in2 => \N__11939\,
            in3 => \N__11912\,
            lcout => \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIKIU51Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FSM_TEST_inst_RAPIDA.current_state_1_rep2_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__11493\,
            in1 => \N__11671\,
            in2 => \N__11749\,
            in3 => \N__11656\,
            lcout => \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10838\,
            ce => 'H',
            sr => \N__10619\
        );

    \FSM_TEST_inst_RAPIDA.current_state_1_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__11670\,
            in1 => \N__11655\,
            in2 => \N__10967\,
            in3 => \N__11494\,
            lcout => \FSM_TEST_inst_RAPIDA.current_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10838\,
            ce => 'H',
            sr => \N__10619\
        );

    \config_register_latched_dec_inst.STATCNF_1_RNIRDN51_0_0_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10454\,
            lcout => \STATCNF_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
