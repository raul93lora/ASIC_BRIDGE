/*
* Raul Lora Rivera
*
* ASIC BRIDGE TOP.v
*
* This module first send to the ASIC analog part the STATCNF and DYNCNF at 2MHz and then at 1MHz
* These frequencies are variable through the DELAY parameters in modules switch_clk_2MHz and switch_clk_1MHz
*
*/
module ASIC_bridge_top(
	CLK,		
	RST_N,
	clk_output,					// Final clock output for Analog ASIC
	static_conf_ear,				// Static configuration register
	dynamic_conf,					// Dynamic configuration register
	mosi_output,					// MOSI signal for Analog ASIC
	sel_output,					// SEL signal for Analog ASIC
	miso_input,					// MISO signal for Analog ASIC
	//s15,						// To test in GPIO the STATCNF or DYNCNF bits				
	//s14,						// To test in GPIO the STATCNF or DYNCNF bits						
	//s13,						// To test in GPIO the STATCNF or DYNCNF bits						
	//s12,						// To test in GPIO the STATCNF or DYNCNF bits
	flag_dyn,
	flag_stat,						
	xor_out_dyn,					// Error for dynamic reg
	xor_out_stat,					// Error for static reg
	start_ASIC_config,				// Input signal to start ASIC config 
	end_config
);

	// Parameters definition
	parameter SIZESRSTAT = 88; 			// Static shift register length 
	parameter SIZESRDYN = 16; 			// Dynamic shift register length
	parameter SIZEADDRMUX = 7;

	// Ports definition
	input wire CLK;
	input wire RST_N;
	input wire miso_input;
	input wire flag_dyn;
	input wire flag_stat;
	input wire [SIZESRSTAT-1:0] static_conf_ear;
	input wire [SIZESRDYN-1:0] dynamic_conf;
	input wire start_ASIC_config;
	output wire clk_output;
	output wire mosi_output;
	output wire sel_output;
	//output wire s15;
	//output wire s14;
	//output wire s13;
	//output wire s12;
	output wire xor_out_dyn;			// Error detection y DYNCNF
	output wire xor_out_stat;			// Error detection y STATCNF
	output wire end_config;

	// Connections
	wire clk_continuous_1MHz;
	wire clk_continuous_2MHz;
	wire clk_out_1MHz;
	wire clk_out_2MHz;
	wire mosi;
	wire mosi_1MHz;
	wire mosi_2MHz;
	wire aux_selection;
	wire aux_selection_1MHz;
	wire aux_selection_2MHz;
	wire clk_output_aux;
	wire mosi_output_aux;
	wire sel_output_aux;
	wire signal_sdo;		
	wire [SIZESRDYN-1:0] DYNLATCH;
	wire [SIZESRSTAT-1:0] STATLATCH;  
	wire [SIZESRDYN-1:0] DYNCNF;
	wire [SIZESRSTAT-1:0] STATCNF;

	// Instantiate frequency divider to generate a continuous 2MHz clock (Fin=16MHz, Fout=2MHz, DIV=8)
	freq_div #(.DIVISOR(8)) divisor_inst (
		.clk_in(CLK),
		.RST_N(RST_N),
		.clk_out(clk_continuous_2MHz)
	);

	// Instantiate switch_clk_2Mhz to switch on/off the 2MHz clock
	switch_clk_write2MHz #(
		.DELAY_CYCLES(8)
    	) switch_clk_write2MHz_STATIC_inst(
		.CLK(CLK),					
		.clk_continuous_2MHz(clk_continuous_2MHz),		
		.CLK_ON_OFF(clk_out_2MHz),					
		.RST_N(RST_N),
		.dynamic_conf(dynamic_conf),
		.static_conf_ear(static_conf_ear),
		.SEL(aux_selection_2MHz),
		.flag_dyn(flag_dyn),
		.flag_stat(flag_stat),
		.end_config(end_config),
		.MOSI(mosi_2MHz),
		.start_ASIC_config(start_ASIC_config)
	);

	// Select between writing at 2MHz or 1MHz
	assign clk_output = clk_out_2MHz;
	assign mosi_output = mosi_2MHz;
	assign sel_output = aux_selection_2MHz;
	//assign s14 = aux_selection_1MHz;
	//assign s13 = aux_selection;

	// Aux signals to choose between 1MHz or 2MHz clock frequencies
	assign clk_output_aux = clk_out_2MHz;
	assign mosi_output_aux = mosi_2MHz;
	assign sel_output_aux = aux_selection_2MHz;

	// Erandel analog chip emulator RTL module (to check that the response from the other FPGA is the same that was sent there)
	config_register_latched_dec config_register_latched_dec_inst(
		.CLK(clk_output_aux), 
		.RST_N(RST_N), 
		.SEL(sel_output_aux), 
		//.SDI(miso_input), 
		.SDI(mosi_output_aux),      				// Simulation and test in the same hardware platform
		.SDO(signal_sdo), 
		.STATCNF(STATCNF), 
		.DYNCNF(DYNCNF), 
		.AMUXSEL(), 
		.STG2_EN(), 
		.STG1_EN(), 
		.ref_elec_en()
	);

	// Error detection for dynamic register (XOR-based detection)
	xor_n_bits #(.N(16)) xor_instance_dyn (
		.a(dynamic_conf),
		.b(DYNCNF),
		.result(xor_out_dyn)
	);

	// Error detection for static register (XOR-based detection)
	xor_n_bits #(.N(88)) xor_instance_stat (
		.a(static_conf_ear),
		.b(STATCNF),
		.result(xor_out_stat)
	);

/*
	// Assignments for output to test correct values for DYNCNF and STATCNF	
	//assign s15 = DYNCNF[7];
	assign s14 = DYNCNF[10];
	assign s13 = DYNCNF[9];
	assign s12 = DYNCNF[8];

	assign s15 = STATCNF[3];
	assign s14 = STATCNF[2];
	assign s13 = STATCNF[1];
	assign s12 = STATCNF[0];
*/


endmodule























