// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 10 2025 16:58:15

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    xor_out_stat,
    mosi_output,
    miso_input,
    xor_out_dyn,
    sel_output,
    s14,
    s12,
    clk_output,
    CLK,
    s13,
    RST_N);

    output xor_out_stat;
    output mosi_output;
    input miso_input;
    output xor_out_dyn;
    output sel_output;
    output s14;
    output s12;
    output clk_output;
    input CLK;
    output s13;
    input RST_N;

    wire N__12279;
    wire N__12278;
    wire N__12277;
    wire N__12270;
    wire N__12269;
    wire N__12268;
    wire N__12261;
    wire N__12260;
    wire N__12259;
    wire N__12252;
    wire N__12251;
    wire N__12250;
    wire N__12243;
    wire N__12242;
    wire N__12241;
    wire N__12234;
    wire N__12233;
    wire N__12232;
    wire N__12225;
    wire N__12224;
    wire N__12223;
    wire N__12216;
    wire N__12215;
    wire N__12214;
    wire N__12207;
    wire N__12206;
    wire N__12205;
    wire N__12198;
    wire N__12197;
    wire N__12196;
    wire N__12189;
    wire N__12188;
    wire N__12187;
    wire N__12170;
    wire N__12167;
    wire N__12164;
    wire N__12161;
    wire N__12158;
    wire N__12155;
    wire N__12152;
    wire N__12151;
    wire N__12150;
    wire N__12149;
    wire N__12148;
    wire N__12147;
    wire N__12146;
    wire N__12145;
    wire N__12144;
    wire N__12143;
    wire N__12142;
    wire N__12141;
    wire N__12140;
    wire N__12139;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12097;
    wire N__12096;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12084;
    wire N__12083;
    wire N__12082;
    wire N__12081;
    wire N__12078;
    wire N__12075;
    wire N__12072;
    wire N__12071;
    wire N__12070;
    wire N__12067;
    wire N__12064;
    wire N__12063;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12035;
    wire N__12034;
    wire N__12025;
    wire N__12022;
    wire N__12019;
    wire N__12016;
    wire N__12011;
    wire N__12008;
    wire N__12005;
    wire N__12002;
    wire N__11999;
    wire N__11998;
    wire N__11997;
    wire N__11996;
    wire N__11993;
    wire N__11992;
    wire N__11985;
    wire N__11982;
    wire N__11979;
    wire N__11972;
    wire N__11969;
    wire N__11968;
    wire N__11965;
    wire N__11964;
    wire N__11961;
    wire N__11960;
    wire N__11957;
    wire N__11954;
    wire N__11951;
    wire N__11948;
    wire N__11939;
    wire N__11936;
    wire N__11935;
    wire N__11934;
    wire N__11931;
    wire N__11930;
    wire N__11925;
    wire N__11922;
    wire N__11919;
    wire N__11912;
    wire N__11911;
    wire N__11910;
    wire N__11909;
    wire N__11908;
    wire N__11905;
    wire N__11902;
    wire N__11895;
    wire N__11892;
    wire N__11885;
    wire N__11882;
    wire N__11879;
    wire N__11876;
    wire N__11873;
    wire N__11872;
    wire N__11871;
    wire N__11870;
    wire N__11869;
    wire N__11868;
    wire N__11867;
    wire N__11866;
    wire N__11865;
    wire N__11864;
    wire N__11863;
    wire N__11862;
    wire N__11861;
    wire N__11854;
    wire N__11853;
    wire N__11852;
    wire N__11851;
    wire N__11848;
    wire N__11847;
    wire N__11836;
    wire N__11835;
    wire N__11834;
    wire N__11833;
    wire N__11832;
    wire N__11831;
    wire N__11830;
    wire N__11829;
    wire N__11828;
    wire N__11827;
    wire N__11826;
    wire N__11825;
    wire N__11824;
    wire N__11821;
    wire N__11818;
    wire N__11813;
    wire N__11812;
    wire N__11811;
    wire N__11810;
    wire N__11807;
    wire N__11802;
    wire N__11795;
    wire N__11792;
    wire N__11781;
    wire N__11772;
    wire N__11765;
    wire N__11760;
    wire N__11757;
    wire N__11750;
    wire N__11749;
    wire N__11744;
    wire N__11741;
    wire N__11736;
    wire N__11731;
    wire N__11724;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11712;
    wire N__11707;
    wire N__11704;
    wire N__11701;
    wire N__11690;
    wire N__11689;
    wire N__11686;
    wire N__11685;
    wire N__11684;
    wire N__11675;
    wire N__11672;
    wire N__11671;
    wire N__11670;
    wire N__11667;
    wire N__11662;
    wire N__11657;
    wire N__11656;
    wire N__11655;
    wire N__11652;
    wire N__11651;
    wire N__11650;
    wire N__11649;
    wire N__11646;
    wire N__11643;
    wire N__11642;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11625;
    wire N__11624;
    wire N__11623;
    wire N__11622;
    wire N__11621;
    wire N__11620;
    wire N__11619;
    wire N__11618;
    wire N__11617;
    wire N__11616;
    wire N__11615;
    wire N__11614;
    wire N__11613;
    wire N__11610;
    wire N__11603;
    wire N__11600;
    wire N__11599;
    wire N__11598;
    wire N__11595;
    wire N__11584;
    wire N__11581;
    wire N__11578;
    wire N__11567;
    wire N__11562;
    wire N__11559;
    wire N__11556;
    wire N__11553;
    wire N__11534;
    wire N__11533;
    wire N__11532;
    wire N__11531;
    wire N__11530;
    wire N__11529;
    wire N__11528;
    wire N__11527;
    wire N__11526;
    wire N__11525;
    wire N__11524;
    wire N__11523;
    wire N__11522;
    wire N__11521;
    wire N__11520;
    wire N__11519;
    wire N__11518;
    wire N__11517;
    wire N__11516;
    wire N__11515;
    wire N__11514;
    wire N__11513;
    wire N__11512;
    wire N__11511;
    wire N__11510;
    wire N__11509;
    wire N__11508;
    wire N__11507;
    wire N__11506;
    wire N__11505;
    wire N__11504;
    wire N__11503;
    wire N__11502;
    wire N__11501;
    wire N__11500;
    wire N__11499;
    wire N__11498;
    wire N__11497;
    wire N__11496;
    wire N__11495;
    wire N__11494;
    wire N__11493;
    wire N__11490;
    wire N__11489;
    wire N__11488;
    wire N__11487;
    wire N__11486;
    wire N__11485;
    wire N__11484;
    wire N__11483;
    wire N__11482;
    wire N__11481;
    wire N__11480;
    wire N__11479;
    wire N__11478;
    wire N__11477;
    wire N__11476;
    wire N__11475;
    wire N__11474;
    wire N__11473;
    wire N__11472;
    wire N__11471;
    wire N__11470;
    wire N__11469;
    wire N__11468;
    wire N__11467;
    wire N__11466;
    wire N__11465;
    wire N__11464;
    wire N__11463;
    wire N__11462;
    wire N__11461;
    wire N__11460;
    wire N__11459;
    wire N__11458;
    wire N__11457;
    wire N__11456;
    wire N__11455;
    wire N__11454;
    wire N__11439;
    wire N__11426;
    wire N__11409;
    wire N__11402;
    wire N__11385;
    wire N__11370;
    wire N__11369;
    wire N__11368;
    wire N__11367;
    wire N__11366;
    wire N__11361;
    wire N__11358;
    wire N__11343;
    wire N__11330;
    wire N__11323;
    wire N__11308;
    wire N__11305;
    wire N__11296;
    wire N__11291;
    wire N__11288;
    wire N__11287;
    wire N__11286;
    wire N__11285;
    wire N__11284;
    wire N__11283;
    wire N__11282;
    wire N__11281;
    wire N__11280;
    wire N__11279;
    wire N__11278;
    wire N__11277;
    wire N__11276;
    wire N__11275;
    wire N__11274;
    wire N__11273;
    wire N__11272;
    wire N__11271;
    wire N__11270;
    wire N__11269;
    wire N__11268;
    wire N__11267;
    wire N__11266;
    wire N__11265;
    wire N__11264;
    wire N__11263;
    wire N__11262;
    wire N__11261;
    wire N__11260;
    wire N__11259;
    wire N__11258;
    wire N__11257;
    wire N__11256;
    wire N__11255;
    wire N__11254;
    wire N__11243;
    wire N__11230;
    wire N__11221;
    wire N__11220;
    wire N__11219;
    wire N__11214;
    wire N__11199;
    wire N__11196;
    wire N__11195;
    wire N__11194;
    wire N__11193;
    wire N__11188;
    wire N__11173;
    wire N__11158;
    wire N__11153;
    wire N__11150;
    wire N__11149;
    wire N__11148;
    wire N__11147;
    wire N__11140;
    wire N__11125;
    wire N__11114;
    wire N__11107;
    wire N__11104;
    wire N__11101;
    wire N__11094;
    wire N__11087;
    wire N__11078;
    wire N__11075;
    wire N__11068;
    wire N__11045;
    wire N__11044;
    wire N__11043;
    wire N__11042;
    wire N__11041;
    wire N__11040;
    wire N__11039;
    wire N__11034;
    wire N__11033;
    wire N__11032;
    wire N__11031;
    wire N__11030;
    wire N__11029;
    wire N__11028;
    wire N__11027;
    wire N__11026;
    wire N__11025;
    wire N__11024;
    wire N__11023;
    wire N__11022;
    wire N__11011;
    wire N__11008;
    wire N__11005;
    wire N__11004;
    wire N__11003;
    wire N__11002;
    wire N__11001;
    wire N__11000;
    wire N__10999;
    wire N__10996;
    wire N__10989;
    wire N__10982;
    wire N__10973;
    wire N__10972;
    wire N__10971;
    wire N__10970;
    wire N__10969;
    wire N__10968;
    wire N__10967;
    wire N__10964;
    wire N__10959;
    wire N__10952;
    wire N__10945;
    wire N__10944;
    wire N__10943;
    wire N__10934;
    wire N__10923;
    wire N__10920;
    wire N__10911;
    wire N__10906;
    wire N__10901;
    wire N__10898;
    wire N__10889;
    wire N__10888;
    wire N__10887;
    wire N__10886;
    wire N__10885;
    wire N__10884;
    wire N__10883;
    wire N__10882;
    wire N__10881;
    wire N__10880;
    wire N__10879;
    wire N__10878;
    wire N__10877;
    wire N__10876;
    wire N__10875;
    wire N__10874;
    wire N__10873;
    wire N__10872;
    wire N__10871;
    wire N__10870;
    wire N__10869;
    wire N__10868;
    wire N__10867;
    wire N__10866;
    wire N__10865;
    wire N__10864;
    wire N__10863;
    wire N__10862;
    wire N__10861;
    wire N__10860;
    wire N__10859;
    wire N__10858;
    wire N__10857;
    wire N__10856;
    wire N__10855;
    wire N__10854;
    wire N__10853;
    wire N__10852;
    wire N__10851;
    wire N__10850;
    wire N__10849;
    wire N__10848;
    wire N__10847;
    wire N__10846;
    wire N__10845;
    wire N__10844;
    wire N__10843;
    wire N__10842;
    wire N__10841;
    wire N__10840;
    wire N__10839;
    wire N__10838;
    wire N__10837;
    wire N__10836;
    wire N__10835;
    wire N__10834;
    wire N__10833;
    wire N__10832;
    wire N__10831;
    wire N__10830;
    wire N__10829;
    wire N__10828;
    wire N__10827;
    wire N__10826;
    wire N__10825;
    wire N__10824;
    wire N__10823;
    wire N__10822;
    wire N__10821;
    wire N__10820;
    wire N__10819;
    wire N__10676;
    wire N__10673;
    wire N__10672;
    wire N__10671;
    wire N__10670;
    wire N__10669;
    wire N__10668;
    wire N__10667;
    wire N__10666;
    wire N__10665;
    wire N__10664;
    wire N__10663;
    wire N__10662;
    wire N__10661;
    wire N__10660;
    wire N__10659;
    wire N__10658;
    wire N__10657;
    wire N__10656;
    wire N__10655;
    wire N__10654;
    wire N__10653;
    wire N__10652;
    wire N__10651;
    wire N__10650;
    wire N__10649;
    wire N__10648;
    wire N__10647;
    wire N__10646;
    wire N__10645;
    wire N__10644;
    wire N__10643;
    wire N__10642;
    wire N__10641;
    wire N__10640;
    wire N__10639;
    wire N__10638;
    wire N__10637;
    wire N__10636;
    wire N__10635;
    wire N__10634;
    wire N__10633;
    wire N__10632;
    wire N__10631;
    wire N__10630;
    wire N__10629;
    wire N__10628;
    wire N__10627;
    wire N__10626;
    wire N__10625;
    wire N__10624;
    wire N__10623;
    wire N__10622;
    wire N__10621;
    wire N__10620;
    wire N__10619;
    wire N__10618;
    wire N__10617;
    wire N__10616;
    wire N__10615;
    wire N__10614;
    wire N__10613;
    wire N__10612;
    wire N__10611;
    wire N__10610;
    wire N__10609;
    wire N__10608;
    wire N__10607;
    wire N__10606;
    wire N__10605;
    wire N__10604;
    wire N__10603;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10342;
    wire N__10341;
    wire N__10340;
    wire N__10339;
    wire N__10338;
    wire N__10337;
    wire N__10336;
    wire N__10335;
    wire N__10334;
    wire N__10333;
    wire N__10332;
    wire N__10331;
    wire N__10330;
    wire N__10329;
    wire N__10328;
    wire N__10327;
    wire N__10326;
    wire N__10325;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10314;
    wire N__10313;
    wire N__10312;
    wire N__10311;
    wire N__10310;
    wire N__10309;
    wire N__10308;
    wire N__10307;
    wire N__10306;
    wire N__10291;
    wire N__10282;
    wire N__10279;
    wire N__10272;
    wire N__10267;
    wire N__10260;
    wire N__10259;
    wire N__10258;
    wire N__10255;
    wire N__10252;
    wire N__10249;
    wire N__10246;
    wire N__10245;
    wire N__10244;
    wire N__10243;
    wire N__10232;
    wire N__10227;
    wire N__10218;
    wire N__10215;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10188;
    wire N__10181;
    wire N__10178;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10153;
    wire N__10150;
    wire N__10149;
    wire N__10146;
    wire N__10143;
    wire N__10140;
    wire N__10137;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10105;
    wire N__10102;
    wire N__10099;
    wire N__10098;
    wire N__10095;
    wire N__10094;
    wire N__10089;
    wire N__10088;
    wire N__10087;
    wire N__10086;
    wire N__10085;
    wire N__10084;
    wire N__10083;
    wire N__10082;
    wire N__10081;
    wire N__10080;
    wire N__10079;
    wire N__10078;
    wire N__10075;
    wire N__10074;
    wire N__10073;
    wire N__10072;
    wire N__10071;
    wire N__10070;
    wire N__10069;
    wire N__10068;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10050;
    wire N__10047;
    wire N__10042;
    wire N__10035;
    wire N__10032;
    wire N__10021;
    wire N__10014;
    wire N__10011;
    wire N__10008;
    wire N__9999;
    wire N__9996;
    wire N__9991;
    wire N__9984;
    wire N__9977;
    wire N__9974;
    wire N__9973;
    wire N__9972;
    wire N__9971;
    wire N__9970;
    wire N__9967;
    wire N__9964;
    wire N__9961;
    wire N__9956;
    wire N__9951;
    wire N__9948;
    wire N__9941;
    wire N__9940;
    wire N__9937;
    wire N__9936;
    wire N__9933;
    wire N__9932;
    wire N__9931;
    wire N__9928;
    wire N__9925;
    wire N__9918;
    wire N__9911;
    wire N__9910;
    wire N__9909;
    wire N__9906;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9881;
    wire N__9880;
    wire N__9879;
    wire N__9878;
    wire N__9877;
    wire N__9874;
    wire N__9873;
    wire N__9866;
    wire N__9863;
    wire N__9860;
    wire N__9857;
    wire N__9854;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9809;
    wire N__9806;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9788;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9653;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9608;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9593;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9581;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9562;
    wire N__9557;
    wire N__9554;
    wire N__9553;
    wire N__9548;
    wire N__9545;
    wire N__9544;
    wire N__9539;
    wire N__9536;
    wire N__9535;
    wire N__9532;
    wire N__9529;
    wire N__9528;
    wire N__9527;
    wire N__9522;
    wire N__9517;
    wire N__9514;
    wire N__9509;
    wire N__9506;
    wire N__9505;
    wire N__9500;
    wire N__9499;
    wire N__9498;
    wire N__9495;
    wire N__9492;
    wire N__9489;
    wire N__9486;
    wire N__9479;
    wire N__9478;
    wire N__9475;
    wire N__9472;
    wire N__9469;
    wire N__9466;
    wire N__9463;
    wire N__9460;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9424;
    wire N__9421;
    wire N__9420;
    wire N__9419;
    wire N__9418;
    wire N__9415;
    wire N__9414;
    wire N__9413;
    wire N__9412;
    wire N__9411;
    wire N__9408;
    wire N__9405;
    wire N__9394;
    wire N__9391;
    wire N__9388;
    wire N__9387;
    wire N__9382;
    wire N__9377;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9343;
    wire N__9340;
    wire N__9337;
    wire N__9332;
    wire N__9331;
    wire N__9326;
    wire N__9323;
    wire N__9322;
    wire N__9317;
    wire N__9314;
    wire N__9313;
    wire N__9310;
    wire N__9307;
    wire N__9302;
    wire N__9301;
    wire N__9296;
    wire N__9293;
    wire N__9292;
    wire N__9291;
    wire N__9290;
    wire N__9289;
    wire N__9288;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9270;
    wire N__9265;
    wire N__9260;
    wire N__9259;
    wire N__9256;
    wire N__9255;
    wire N__9254;
    wire N__9251;
    wire N__9250;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9240;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9221;
    wire N__9216;
    wire N__9213;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9196;
    wire N__9193;
    wire N__9192;
    wire N__9189;
    wire N__9186;
    wire N__9183;
    wire N__9182;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9164;
    wire N__9163;
    wire N__9162;
    wire N__9161;
    wire N__9160;
    wire N__9153;
    wire N__9148;
    wire N__9145;
    wire N__9140;
    wire N__9139;
    wire N__9136;
    wire N__9135;
    wire N__9134;
    wire N__9131;
    wire N__9130;
    wire N__9129;
    wire N__9122;
    wire N__9115;
    wire N__9110;
    wire N__9109;
    wire N__9108;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9091;
    wire N__9086;
    wire N__9085;
    wire N__9082;
    wire N__9081;
    wire N__9078;
    wire N__9075;
    wire N__9072;
    wire N__9069;
    wire N__9062;
    wire N__9061;
    wire N__9060;
    wire N__9057;
    wire N__9052;
    wire N__9051;
    wire N__9050;
    wire N__9049;
    wire N__9048;
    wire N__9047;
    wire N__9046;
    wire N__9045;
    wire N__9044;
    wire N__9043;
    wire N__9042;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9030;
    wire N__9029;
    wire N__9028;
    wire N__9027;
    wire N__9026;
    wire N__9025;
    wire N__9024;
    wire N__9023;
    wire N__9022;
    wire N__9021;
    wire N__9020;
    wire N__9019;
    wire N__9018;
    wire N__9017;
    wire N__9016;
    wire N__9015;
    wire N__9014;
    wire N__9013;
    wire N__9012;
    wire N__9011;
    wire N__9010;
    wire N__9009;
    wire N__9008;
    wire N__9007;
    wire N__9006;
    wire N__9005;
    wire N__9004;
    wire N__9003;
    wire N__9002;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8988;
    wire N__8987;
    wire N__8986;
    wire N__8985;
    wire N__8984;
    wire N__8983;
    wire N__8982;
    wire N__8981;
    wire N__8980;
    wire N__8979;
    wire N__8978;
    wire N__8977;
    wire N__8976;
    wire N__8975;
    wire N__8974;
    wire N__8973;
    wire N__8972;
    wire N__8971;
    wire N__8970;
    wire N__8969;
    wire N__8968;
    wire N__8967;
    wire N__8966;
    wire N__8965;
    wire N__8964;
    wire N__8963;
    wire N__8962;
    wire N__8961;
    wire N__8960;
    wire N__8959;
    wire N__8958;
    wire N__8957;
    wire N__8956;
    wire N__8955;
    wire N__8954;
    wire N__8953;
    wire N__8952;
    wire N__8951;
    wire N__8950;
    wire N__8947;
    wire N__8942;
    wire N__8941;
    wire N__8940;
    wire N__8939;
    wire N__8938;
    wire N__8937;
    wire N__8936;
    wire N__8935;
    wire N__8934;
    wire N__8933;
    wire N__8932;
    wire N__8931;
    wire N__8930;
    wire N__8927;
    wire N__8920;
    wire N__8909;
    wire N__8898;
    wire N__8883;
    wire N__8880;
    wire N__8863;
    wire N__8858;
    wire N__8857;
    wire N__8856;
    wire N__8855;
    wire N__8854;
    wire N__8851;
    wire N__8848;
    wire N__8845;
    wire N__8834;
    wire N__8827;
    wire N__8824;
    wire N__8817;
    wire N__8804;
    wire N__8789;
    wire N__8778;
    wire N__8769;
    wire N__8768;
    wire N__8765;
    wire N__8756;
    wire N__8751;
    wire N__8742;
    wire N__8725;
    wire N__8724;
    wire N__8723;
    wire N__8722;
    wire N__8721;
    wire N__8720;
    wire N__8719;
    wire N__8718;
    wire N__8717;
    wire N__8716;
    wire N__8715;
    wire N__8714;
    wire N__8713;
    wire N__8712;
    wire N__8711;
    wire N__8710;
    wire N__8709;
    wire N__8698;
    wire N__8695;
    wire N__8690;
    wire N__8681;
    wire N__8670;
    wire N__8657;
    wire N__8654;
    wire N__8653;
    wire N__8652;
    wire N__8651;
    wire N__8650;
    wire N__8645;
    wire N__8640;
    wire N__8637;
    wire N__8626;
    wire N__8611;
    wire N__8604;
    wire N__8601;
    wire N__8592;
    wire N__8585;
    wire N__8576;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8536;
    wire N__8535;
    wire N__8534;
    wire N__8533;
    wire N__8530;
    wire N__8527;
    wire N__8520;
    wire N__8513;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8503;
    wire N__8498;
    wire N__8497;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8486;
    wire N__8483;
    wire N__8478;
    wire N__8475;
    wire N__8468;
    wire N__8467;
    wire N__8464;
    wire N__8463;
    wire N__8462;
    wire N__8457;
    wire N__8456;
    wire N__8455;
    wire N__8454;
    wire N__8451;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8434;
    wire N__8433;
    wire N__8432;
    wire N__8429;
    wire N__8420;
    wire N__8415;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8383;
    wire N__8380;
    wire N__8375;
    wire N__8372;
    wire N__8369;
    wire N__8366;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8354;
    wire N__8353;
    wire N__8352;
    wire N__8351;
    wire N__8350;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8327;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8309;
    wire N__8306;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8273;
    wire N__8270;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8233;
    wire N__8232;
    wire N__8229;
    wire N__8226;
    wire N__8223;
    wire N__8218;
    wire N__8215;
    wire N__8210;
    wire N__8207;
    wire N__8204;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8191;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8179;
    wire N__8176;
    wire N__8175;
    wire N__8172;
    wire N__8169;
    wire N__8166;
    wire N__8163;
    wire N__8156;
    wire N__8155;
    wire N__8150;
    wire N__8147;
    wire N__8144;
    wire N__8141;
    wire N__8138;
    wire N__8135;
    wire N__8132;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8124;
    wire N__8123;
    wire N__8118;
    wire N__8113;
    wire N__8110;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8068;
    wire N__8063;
    wire N__8062;
    wire N__8061;
    wire N__8058;
    wire N__8053;
    wire N__8050;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8033;
    wire N__8030;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7990;
    wire N__7985;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7939;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7931;
    wire N__7930;
    wire N__7929;
    wire N__7928;
    wire N__7927;
    wire N__7926;
    wire N__7925;
    wire N__7924;
    wire N__7923;
    wire N__7922;
    wire N__7921;
    wire N__7920;
    wire N__7919;
    wire N__7918;
    wire N__7917;
    wire N__7916;
    wire N__7915;
    wire N__7914;
    wire N__7913;
    wire N__7910;
    wire N__7909;
    wire N__7908;
    wire N__7907;
    wire N__7906;
    wire N__7905;
    wire N__7904;
    wire N__7903;
    wire N__7902;
    wire N__7901;
    wire N__7900;
    wire N__7899;
    wire N__7892;
    wire N__7889;
    wire N__7888;
    wire N__7887;
    wire N__7886;
    wire N__7885;
    wire N__7882;
    wire N__7881;
    wire N__7880;
    wire N__7879;
    wire N__7878;
    wire N__7877;
    wire N__7876;
    wire N__7875;
    wire N__7872;
    wire N__7869;
    wire N__7866;
    wire N__7865;
    wire N__7864;
    wire N__7863;
    wire N__7860;
    wire N__7859;
    wire N__7858;
    wire N__7855;
    wire N__7852;
    wire N__7851;
    wire N__7850;
    wire N__7849;
    wire N__7848;
    wire N__7845;
    wire N__7842;
    wire N__7841;
    wire N__7838;
    wire N__7837;
    wire N__7836;
    wire N__7835;
    wire N__7834;
    wire N__7833;
    wire N__7832;
    wire N__7831;
    wire N__7830;
    wire N__7829;
    wire N__7828;
    wire N__7827;
    wire N__7824;
    wire N__7821;
    wire N__7818;
    wire N__7815;
    wire N__7814;
    wire N__7813;
    wire N__7812;
    wire N__7811;
    wire N__7808;
    wire N__7807;
    wire N__7804;
    wire N__7801;
    wire N__7800;
    wire N__7799;
    wire N__7798;
    wire N__7797;
    wire N__7796;
    wire N__7791;
    wire N__7786;
    wire N__7785;
    wire N__7782;
    wire N__7781;
    wire N__7778;
    wire N__7775;
    wire N__7774;
    wire N__7773;
    wire N__7770;
    wire N__7767;
    wire N__7766;
    wire N__7763;
    wire N__7762;
    wire N__7761;
    wire N__7758;
    wire N__7757;
    wire N__7754;
    wire N__7753;
    wire N__7752;
    wire N__7749;
    wire N__7746;
    wire N__7743;
    wire N__7736;
    wire N__7733;
    wire N__7722;
    wire N__7707;
    wire N__7700;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7671;
    wire N__7670;
    wire N__7669;
    wire N__7668;
    wire N__7667;
    wire N__7666;
    wire N__7665;
    wire N__7664;
    wire N__7663;
    wire N__7654;
    wire N__7645;
    wire N__7644;
    wire N__7641;
    wire N__7640;
    wire N__7639;
    wire N__7638;
    wire N__7635;
    wire N__7632;
    wire N__7621;
    wire N__7620;
    wire N__7617;
    wire N__7614;
    wire N__7609;
    wire N__7602;
    wire N__7593;
    wire N__7588;
    wire N__7573;
    wire N__7572;
    wire N__7571;
    wire N__7570;
    wire N__7569;
    wire N__7568;
    wire N__7567;
    wire N__7566;
    wire N__7565;
    wire N__7564;
    wire N__7563;
    wire N__7562;
    wire N__7561;
    wire N__7548;
    wire N__7537;
    wire N__7536;
    wire N__7535;
    wire N__7534;
    wire N__7525;
    wire N__7514;
    wire N__7509;
    wire N__7504;
    wire N__7487;
    wire N__7482;
    wire N__7471;
    wire N__7468;
    wire N__7463;
    wire N__7460;
    wire N__7459;
    wire N__7458;
    wire N__7457;
    wire N__7454;
    wire N__7447;
    wire N__7444;
    wire N__7439;
    wire N__7432;
    wire N__7427;
    wire N__7420;
    wire N__7411;
    wire N__7406;
    wire N__7399;
    wire N__7392;
    wire N__7383;
    wire N__7376;
    wire N__7369;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7333;
    wire N__7332;
    wire N__7331;
    wire N__7330;
    wire N__7329;
    wire N__7328;
    wire N__7327;
    wire N__7326;
    wire N__7325;
    wire N__7324;
    wire N__7323;
    wire N__7322;
    wire N__7321;
    wire N__7320;
    wire N__7319;
    wire N__7318;
    wire N__7317;
    wire N__7316;
    wire N__7315;
    wire N__7314;
    wire N__7313;
    wire N__7312;
    wire N__7311;
    wire N__7310;
    wire N__7259;
    wire N__7256;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7244;
    wire N__7241;
    wire N__7240;
    wire N__7239;
    wire N__7238;
    wire N__7235;
    wire N__7228;
    wire N__7227;
    wire N__7226;
    wire N__7225;
    wire N__7222;
    wire N__7219;
    wire N__7212;
    wire N__7211;
    wire N__7210;
    wire N__7209;
    wire N__7208;
    wire N__7205;
    wire N__7200;
    wire N__7191;
    wire N__7184;
    wire N__7181;
    wire N__7178;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7166;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7136;
    wire N__7133;
    wire N__7130;
    wire N__7127;
    wire N__7124;
    wire N__7121;
    wire N__7118;
    wire N__7115;
    wire N__7112;
    wire N__7109;
    wire N__7106;
    wire N__7103;
    wire N__7100;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7073;
    wire N__7070;
    wire N__7067;
    wire N__7064;
    wire N__7061;
    wire N__7058;
    wire N__7055;
    wire N__7052;
    wire N__7049;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7021;
    wire N__7018;
    wire N__7017;
    wire N__7014;
    wire N__7011;
    wire N__7008;
    wire N__7005;
    wire N__7002;
    wire N__6999;
    wire N__6992;
    wire N__6989;
    wire N__6986;
    wire N__6985;
    wire N__6984;
    wire N__6983;
    wire N__6980;
    wire N__6977;
    wire N__6972;
    wire N__6965;
    wire N__6962;
    wire N__6959;
    wire N__6956;
    wire N__6953;
    wire N__6950;
    wire N__6947;
    wire N__6944;
    wire N__6943;
    wire N__6942;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6928;
    wire N__6925;
    wire N__6920;
    wire N__6917;
    wire N__6916;
    wire N__6913;
    wire N__6912;
    wire N__6909;
    wire N__6908;
    wire N__6905;
    wire N__6898;
    wire N__6893;
    wire N__6892;
    wire N__6891;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6866;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6832;
    wire N__6829;
    wire N__6824;
    wire N__6821;
    wire N__6820;
    wire N__6815;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6800;
    wire N__6799;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6755;
    wire N__6752;
    wire N__6749;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6718;
    wire N__6717;
    wire N__6716;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6697;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6659;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6644;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6617;
    wire N__6616;
    wire N__6613;
    wire N__6610;
    wire N__6609;
    wire N__6606;
    wire N__6603;
    wire N__6602;
    wire N__6599;
    wire N__6596;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6557;
    wire N__6554;
    wire N__6551;
    wire N__6548;
    wire N__6545;
    wire N__6542;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6530;
    wire N__6529;
    wire N__6528;
    wire N__6525;
    wire N__6522;
    wire N__6521;
    wire N__6520;
    wire N__6517;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6501;
    wire N__6498;
    wire N__6491;
    wire N__6488;
    wire N__6487;
    wire N__6486;
    wire N__6485;
    wire N__6484;
    wire N__6475;
    wire N__6472;
    wire N__6467;
    wire N__6464;
    wire N__6461;
    wire N__6460;
    wire N__6459;
    wire N__6456;
    wire N__6453;
    wire N__6450;
    wire N__6445;
    wire N__6440;
    wire N__6439;
    wire N__6438;
    wire N__6435;
    wire N__6434;
    wire N__6431;
    wire N__6424;
    wire N__6419;
    wire N__6418;
    wire N__6417;
    wire N__6412;
    wire N__6409;
    wire N__6404;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6380;
    wire N__6377;
    wire N__6374;
    wire N__6371;
    wire N__6368;
    wire N__6365;
    wire N__6362;
    wire N__6359;
    wire N__6356;
    wire N__6353;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6326;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6316;
    wire N__6315;
    wire N__6314;
    wire N__6311;
    wire N__6304;
    wire N__6299;
    wire N__6298;
    wire N__6295;
    wire N__6294;
    wire N__6293;
    wire N__6290;
    wire N__6283;
    wire N__6278;
    wire N__6277;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6267;
    wire N__6264;
    wire N__6261;
    wire N__6254;
    wire N__6251;
    wire N__6250;
    wire N__6249;
    wire N__6248;
    wire N__6245;
    wire N__6244;
    wire N__6241;
    wire N__6238;
    wire N__6237;
    wire N__6234;
    wire N__6233;
    wire N__6230;
    wire N__6217;
    wire N__6212;
    wire N__6211;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6185;
    wire N__6184;
    wire N__6181;
    wire N__6180;
    wire N__6177;
    wire N__6174;
    wire N__6171;
    wire N__6168;
    wire N__6165;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6131;
    wire N__6128;
    wire N__6125;
    wire N__6124;
    wire N__6123;
    wire N__6118;
    wire N__6115;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6103;
    wire N__6102;
    wire N__6097;
    wire N__6094;
    wire N__6089;
    wire N__6086;
    wire N__6083;
    wire N__6080;
    wire N__6079;
    wire N__6078;
    wire N__6077;
    wire N__6074;
    wire N__6069;
    wire N__6066;
    wire N__6059;
    wire N__6056;
    wire N__6053;
    wire N__6052;
    wire N__6051;
    wire N__6048;
    wire N__6045;
    wire N__6042;
    wire N__6035;
    wire N__6032;
    wire N__6029;
    wire N__6028;
    wire N__6027;
    wire N__6026;
    wire N__6023;
    wire N__6020;
    wire N__6015;
    wire N__6008;
    wire N__6007;
    wire N__6006;
    wire N__6005;
    wire N__6002;
    wire N__5999;
    wire N__5994;
    wire N__5987;
    wire N__5986;
    wire N__5985;
    wire N__5984;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5963;
    wire N__5962;
    wire N__5959;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5942;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5911;
    wire N__5910;
    wire N__5907;
    wire N__5904;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5843;
    wire N__5840;
    wire N__5837;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5825;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5759;
    wire N__5756;
    wire N__5753;
    wire N__5750;
    wire N__5749;
    wire N__5748;
    wire N__5745;
    wire N__5742;
    wire N__5739;
    wire N__5732;
    wire N__5729;
    wire N__5726;
    wire N__5725;
    wire N__5724;
    wire N__5721;
    wire N__5720;
    wire N__5719;
    wire N__5718;
    wire N__5715;
    wire N__5704;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5689;
    wire N__5688;
    wire N__5685;
    wire N__5682;
    wire N__5679;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5656;
    wire N__5655;
    wire N__5654;
    wire N__5645;
    wire N__5644;
    wire N__5643;
    wire N__5642;
    wire N__5641;
    wire N__5638;
    wire N__5629;
    wire N__5624;
    wire N__5623;
    wire N__5622;
    wire N__5619;
    wire N__5616;
    wire N__5613;
    wire N__5606;
    wire N__5605;
    wire N__5604;
    wire N__5601;
    wire N__5598;
    wire N__5595;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5525;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5513;
    wire N__5510;
    wire N__5509;
    wire N__5506;
    wire N__5505;
    wire N__5502;
    wire N__5499;
    wire N__5496;
    wire N__5489;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5467;
    wire N__5466;
    wire N__5465;
    wire N__5460;
    wire N__5455;
    wire N__5450;
    wire N__5449;
    wire N__5446;
    wire N__5445;
    wire N__5442;
    wire N__5437;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5390;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5348;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5336;
    wire N__5333;
    wire N__5330;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5048;
    wire N__5045;
    wire N__5042;
    wire N__5039;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5005;
    wire N__5002;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4940;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire GNDG0;
    wire CLK_c;
    wire VCCG0;
    wire DYNCNF_i_0;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_49 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_38 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_34 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_35 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_36 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_37 ;
    wire \FSM_TEST_inst_slow.CLK_uCZ0 ;
    wire \FSM_TEST_inst_slow.CLK_uC_6c_0_0 ;
    wire \FSM_TEST_inst_slow.CLK_uC_6b_0_0 ;
    wire \FSM_TEST_inst_slow.CLK_uC_2_0_0 ;
    wire \FSM_TEST_inst_slow.CLK_uC_5_0_0 ;
    wire \FSM_TEST_inst_slow.CLK_uC_6_0_0 ;
    wire \FSM_TEST_inst_slow.CLK_uC_6dZ0Z_0 ;
    wire \FSM_TEST_inst_slow.CLK_uC_6eZ0Z_0 ;
    wire \FSM_TEST_inst_slow.CLK_uC_6fZ0Z_0 ;
    wire \FSM_TEST_inst_slow.CLK_uC_3_0_0 ;
    wire \FSM_TEST_inst_slow.CLK_uC_4_0_0 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_16 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_17 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_33 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_48 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_30 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_71 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_31 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_32 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_72 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_41 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_39 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_40 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_12 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_13 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_3 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_2 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_11 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_14 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_4 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_5 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_6 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_7 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_8 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_9 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_10 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_0 ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_1 ;
    wire \FSM_TEST_inst_slow.CLK_uC_6iZ0Z_0 ;
    wire \FSM_TEST_inst_slow.CLK_uC_6jZ0Z_0 ;
    wire \FSM_TEST_inst_slow.CLK_uC_6gZ0Z_0 ;
    wire \FSM_TEST_inst_slow.CLK_uC_6hZ0Z_0 ;
    wire bfn_9_20_0_;
    wire \FSM_TEST_inst_RAPIDA.counter_stat_cry_0 ;
    wire \FSM_TEST_inst_RAPIDA.counter_stat_cry_1 ;
    wire \FSM_TEST_inst_RAPIDA.counter_stat_cry_2 ;
    wire \FSM_TEST_inst_RAPIDA.counter_stat_cry_3 ;
    wire \FSM_TEST_inst_RAPIDA.counter_stat_cry_4 ;
    wire \FSM_TEST_inst_RAPIDA.counter_stat_cry_5 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_15 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_14 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_22 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_20 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_21 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_18 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_19 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_25 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_26 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_29 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_23 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_24 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_27 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_28 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_47 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_73 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_74 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_75 ;
    wire \FSM_TEST_inst_slow.N_134_1_cascade_ ;
    wire \FSM_TEST_inst_slow.bit_sequence_dinZ0Z_15 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_87 ;
    wire \FSM_TEST_inst_slow.G_31_1 ;
    wire \FSM_TEST_inst_slow.counter_statlde_0_cascade_ ;
    wire \FSM_TEST_inst_slow.current_state_RNIR2L81Z0Z_1 ;
    wire bfn_10_18_0_;
    wire \FSM_TEST_inst_slow.counter_idle_cry_0 ;
    wire \FSM_TEST_inst_slow.counter_idle_cry_1 ;
    wire \FSM_TEST_inst_slow.counter_idle_cry_2 ;
    wire \FSM_TEST_inst_slow.counter_idle_cry_3 ;
    wire \FSM_TEST_inst_slow.counter_idle_cry_4 ;
    wire \FSM_TEST_inst_slow.counter_idle_cry_5 ;
    wire \FSM_TEST_inst_slow.counter_idle_cry_6 ;
    wire \FSM_TEST_inst_slow.counter_idle_RNIHR3A2Z0Z_7 ;
    wire \FSM_TEST_inst_slow.counter_idleZ0Z_1 ;
    wire \FSM_TEST_inst_slow.counter_idleZ0Z_2 ;
    wire \FSM_TEST_inst_slow.counter_idleZ0Z_5 ;
    wire \FSM_TEST_inst_slow.counter_idleZ0Z_0 ;
    wire \FSM_TEST_inst_slow.N_109_0 ;
    wire \FSM_TEST_inst_slow.counter_dinZ0Z_0 ;
    wire \FSM_TEST_inst_slow.counter_dinZ1Z_1 ;
    wire \FSM_TEST_inst_slow.N_134_1_i ;
    wire \FSM_TEST_inst_slow.counter_idleZ0Z_4 ;
    wire \FSM_TEST_inst_slow.counter_idleZ0Z_3 ;
    wire \FSM_TEST_inst_RAPIDA.counter_stat_cry_3_THRU_CO ;
    wire \FSM_TEST_inst_RAPIDA.counter_stat_cry_4_THRU_CO ;
    wire \FSM_TEST_inst_RAPIDA.counter_stat_cry_2_THRU_CO ;
    wire \FSM_TEST_inst_RAPIDA.counter_statlde_0_cascade_ ;
    wire \FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2Z0Z_1_cascade_ ;
    wire \FSM_TEST_inst_RAPIDA.counter_statZ0Z_0 ;
    wire \FSM_TEST_inst_RAPIDA.counter_stat_cry_0_THRU_CO ;
    wire \FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2Z0Z_1 ;
    wire \FSM_TEST_inst_RAPIDA.counter_stat_cry_1_THRU_CO ;
    wire \FSM_TEST_inst_RAPIDA.counter_statZ0Z_2 ;
    wire bfn_10_21_0_;
    wire \FSM_TEST_inst_RAPIDA.counter_idle_cry_0 ;
    wire \FSM_TEST_inst_RAPIDA.counter_idle_cry_1 ;
    wire \FSM_TEST_inst_RAPIDA.counter_idle_cry_2 ;
    wire \FSM_TEST_inst_RAPIDA.counter_idle_cry_3 ;
    wire \FSM_TEST_inst_RAPIDA.counter_idle_cry_4 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_13 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_0 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_81 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_46 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_4 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_1 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_2 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_3 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_80 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_42 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_70 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_45 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_76 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_77 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_43 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_44 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_78 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_79 ;
    wire bfn_11_17_0_;
    wire \FSM_TEST_inst_slow.counter_stat_cry_0 ;
    wire \FSM_TEST_inst_slow.counter_stat_cry_1 ;
    wire \FSM_TEST_inst_slow.counter_stat_cry_2 ;
    wire \FSM_TEST_inst_slow.counter_stat_cry_3 ;
    wire \FSM_TEST_inst_slow.counter_stat_cry_4 ;
    wire \FSM_TEST_inst_slow.counter_stat_cry_5 ;
    wire \FSM_TEST_inst_slow.counter_statZ0Z_6 ;
    wire \FSM_TEST_inst_slow.current_state_ns_0_a3_1_4_0_cascade_ ;
    wire \FSM_TEST_inst_slow.current_state_ns_0_a3_1_5_0 ;
    wire \FSM_TEST_inst_slow.counter_statZ0Z_0 ;
    wire \FSM_TEST_inst_slow.counter_stat_cry_1_THRU_CO ;
    wire \FSM_TEST_inst_slow.counter_statZ0Z_2 ;
    wire \FSM_TEST_inst_slow.counter_stat_cry_2_THRU_CO ;
    wire \FSM_TEST_inst_slow.counter_statZ0Z_3 ;
    wire \FSM_TEST_inst_slow.counter_stat_cry_0_THRU_CO ;
    wire \FSM_TEST_inst_slow.counter_statZ0Z_1 ;
    wire \FSM_TEST_inst_slow.counter_stat_cry_3_THRU_CO ;
    wire \FSM_TEST_inst_slow.counter_statZ0Z_4 ;
    wire \FSM_TEST_inst_RAPIDA.counter_statZ0Z_4 ;
    wire \FSM_TEST_inst_RAPIDA.counter_statZ0Z_5 ;
    wire \FSM_TEST_inst_RAPIDA.counter_statZ0Z_1 ;
    wire \FSM_TEST_inst_RAPIDA.counter_idle_cry_0_THRU_CO ;
    wire \FSM_TEST_inst_RAPIDA.N_126_1_i_cascade_ ;
    wire \FSM_TEST_inst_RAPIDA.current_state_d_i_2 ;
    wire \FSM_TEST_inst_slow.counter_idleZ0Z_7 ;
    wire \FSM_TEST_inst_slow.flag_input_regZ0 ;
    wire \FSM_TEST_inst_slow.counter_idleZ0Z_6 ;
    wire \FSM_TEST_inst_slow.current_state_RNO_3Z0Z_0 ;
    wire \FSM_TEST_inst_slow.current_state_RNO_4Z0Z_0_cascade_ ;
    wire \FSM_TEST_inst_slow.current_state_RNO_5Z0Z_0 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_0 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_1 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_2 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_3 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_4 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_5 ;
    wire \FSM_TEST_inst_RAPIDA.counter_idle_cry_3_THRU_CO ;
    wire \FSM_TEST_inst_RAPIDA.flag_input_regZ0 ;
    wire \FSM_TEST_inst_RAPIDA.G_24_0_a4_1_4 ;
    wire \FSM_TEST_inst_RAPIDA.counter_idle_cry_1_THRU_CO ;
    wire \FSM_TEST_inst_RAPIDA.counter_idle_cry_2_THRU_CO ;
    wire \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_4 ;
    wire \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_3 ;
    wire \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_5 ;
    wire \FSM_TEST_inst_RAPIDA.counter_idlelde_2_cascade_ ;
    wire \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1 ;
    wire \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1_cascade_ ;
    wire \FSM_TEST_inst_RAPIDA.N_126_1_i ;
    wire \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_1 ;
    wire \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_2 ;
    wire \FSM_TEST_inst_RAPIDA.counter_idleZ0Z_0 ;
    wire \FSM_TEST_inst_RAPIDA.G_24_0_a4_1_5 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_6 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_19 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_20 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_21 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_22 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_23 ;
    wire CONSTANT_ONE_NET;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_86 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_84 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_85 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_82 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_83 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_12 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_52 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_7 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_8 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_9 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_53 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_10 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_11 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_54 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_55 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_50 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_51 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_5 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_6 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_56 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_69 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_68 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_67 ;
    wire \FSM_TEST_inst_slow.N_108_li_cascade_ ;
    wire \FSM_TEST_inst_slow.current_state_RNIR2L81_0Z0Z_1 ;
    wire \FSM_TEST_inst_slow.current_state_cnv_0_1 ;
    wire \FSM_TEST_inst_slow.N_108_li ;
    wire \FSM_TEST_inst_slow.counter_dinZ0Z_3 ;
    wire \FSM_TEST_inst_slow.counter_dinZ0Z_2 ;
    wire \FSM_TEST_inst_slow.N_106_0 ;
    wire \FSM_TEST_inst_slow.current_state_RNO_8Z0Z_0_cascade_ ;
    wire \FSM_TEST_inst_slow.current_state_RNO_1Z0Z_0 ;
    wire \FSM_TEST_inst_slow.N_134 ;
    wire \FSM_TEST_inst_slow.current_state_RNO_2Z0Z_0_cascade_ ;
    wire s12_c;
    wire \config_register_latched_dec_inst.DYNCNF_1Z0Z_8 ;
    wire \config_register_latched_dec_inst.DYNCNF_1Z0Z_9 ;
    wire s13_c;
    wire \config_register_latched_dec_inst.DYNCNF_1Z0Z_0 ;
    wire \config_register_latched_dec_inst.DYNCNF_0 ;
    wire \FSM_TEST_inst_RAPIDA.counter_din_3_i_0_2_cascade_ ;
    wire \FSM_TEST_inst_RAPIDA.G_24_0_o4_2_cascade_ ;
    wire \FSM_TEST_inst_RAPIDA.G_24_0_a4_0_1 ;
    wire \FSM_TEST_inst_RAPIDA.counter_statZ0Z_6 ;
    wire \FSM_TEST_inst_RAPIDA.counter_statZ0Z_3 ;
    wire \FSM_TEST_inst_RAPIDA.G_24_0_a4_0_5 ;
    wire \FSM_TEST_inst_RAPIDA.N_18_0 ;
    wire \FSM_TEST_inst_RAPIDA.G_24_0_a4_0_6_cascade_ ;
    wire \FSM_TEST_inst_RAPIDA.N_9_1 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_0 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_1 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_4 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_5 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_2 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_3 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_13 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_14 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_18 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_24 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_78 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_77 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_25 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_26 ;
    wire \FSM_TEST_inst_RAPIDA.CLK_uC_3Z0Z_0 ;
    wire \FSM_TEST_inst_RAPIDA.CLK_uC_4Z0Z_0 ;
    wire \FSM_TEST_inst_RAPIDA.CLK_uC_5Z0Z_0 ;
    wire \FSM_TEST_inst_RAPIDA.CLK_uC_6Z0Z_0 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_57 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_60 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_58 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_59 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_61 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_66 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_64 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_65 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_62 ;
    wire \FSM_TEST_inst_slow.current_stateZ0Z_1 ;
    wire \FSM_TEST_inst_slow.bit_sequence_statZ0Z_63 ;
    wire \FSM_TEST_inst_slow.N_374_g ;
    wire counter_RNIFD27_2_cascade_;
    wire N_3_0_cascade_;
    wire N_2_0;
    wire counter_RNISR1F_2;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_15 ;
    wire clk_out_RNI3LEM_cascade_;
    wire \FSM_TEST_inst_RAPIDA.N_100_li_cascade_ ;
    wire \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5DZ0Z1_cascade_ ;
    wire N_378_i;
    wire flag_signal;
    wire mosi_fast;
    wire mosi_slow;
    wire mosi_output_c;
    wire \config_register_latched_dec_inst.DYNCNF_1Z0Z_10 ;
    wire s14_c;
    wire \config_register_latched_dec_inst.N_378_i_i ;
    wire \FSM_TEST_inst_RAPIDA.N_101_0 ;
    wire \config_register_latched_dec_inst.DYNSRZ0Z_10 ;
    wire miso_input_c;
    wire \config_register_latched_dec_inst.DYNSRZ0Z_0 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_10 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_6 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_7 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_8 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_9 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_11 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_12 ;
    wire \FSM_TEST_inst_RAPIDA.current_state_fast_RNI78E11Z0Z_1 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_27 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_28 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_59 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_76 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_54 ;
    wire \FSM_TEST_inst_RAPIDA.CLK_uC_2Z0Z_0 ;
    wire \FSM_TEST_inst_RAPIDA.CLK_uC_6bZ0Z_0 ;
    wire \FSM_TEST_inst_RAPIDA.CLK_uCZ0 ;
    wire \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5DZ0Z1 ;
    wire N_3_0;
    wire N_4_0;
    wire CLK_uC_6c_0;
    wire clk_output_c;
    wire \FSM_TEST_inst_slow.current_state_RNI9C3K2Z0Z_1 ;
    wire \FSM_TEST_inst_slow.current_state_d_i_2 ;
    wire \FSM_TEST_inst_slow.counter_stat_cry_4_THRU_CO ;
    wire \FSM_TEST_inst_slow.counter_statZ0Z_5 ;
    wire \divisor_inst_2.counterZ0Z_1 ;
    wire \divisor_inst_2.counterZ0Z_0 ;
    wire \divisor_inst_2.counterZ0Z_2 ;
    wire \FSM_TEST_inst_RAPIDA.aux_selection_fast_0 ;
    wire \FSM_TEST_inst_slow.current_stateZ1Z_0 ;
    wire counter_RNIFD27_2;
    wire clk_continuous_slow;
    wire \FSM_TEST_inst_slow.aux_selection_slow_0 ;
    wire \FSM_TEST_inst_RAPIDA.current_state_fast_fastZ0Z_1 ;
    wire \FSM_TEST_inst_RAPIDA.current_state_fast_1_repZ0Z1 ;
    wire \FSM_TEST_inst_RAPIDA.current_state_fastZ0Z_1 ;
    wire \FSM_TEST_inst_slow.CLK_uC_6kZ0Z_0 ;
    wire CLK_uC_6l_0;
    wire \config_register_latched_dec_inst.DYNSRZ0Z_3 ;
    wire \config_register_latched_dec_inst.DYNSRZ0Z_4 ;
    wire \config_register_latched_dec_inst.DYNSRZ0Z_1 ;
    wire \config_register_latched_dec_inst.DYNSRZ0Z_2 ;
    wire \config_register_latched_dec_inst.DYNSRZ0Z_7 ;
    wire \config_register_latched_dec_inst.DYNSRZ0Z_5 ;
    wire \config_register_latched_dec_inst.DYNSRZ0Z_6 ;
    wire \config_register_latched_dec_inst.DYNSRZ0Z_8 ;
    wire \config_register_latched_dec_inst.DYNSRZ0Z_9 ;
    wire flag_output_0_ret_RNI1E8NZ0Z2;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_51 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_52 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_53 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_31 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_50 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_29 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_30 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_75 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_60 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_58 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_7 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_8 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_9 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_57 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_79 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_55 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_56 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_83 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_87 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_84 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_85 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_86 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_82 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_65 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_35 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_80 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_81 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_32 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_39 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_46 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_47 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_40 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_48 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_49 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_33 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_34 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_10 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_74 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_13 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_14 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_15 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_16 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_17 ;
    wire \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z1 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_11 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_12 ;
    wire \config_register_latched_dec_inst.STATSRZ0Z_0 ;
    wire \config_register_latched_dec_inst.STATCNF_1Z0Z_0 ;
    wire sel_output_c;
    wire \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_2 ;
    wire \FSM_TEST_inst_RAPIDA.counter_dinZ1Z_1 ;
    wire \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_3 ;
    wire \FSM_TEST_inst_RAPIDA.counter_dinZ0Z_0 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_66 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_67 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_45 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_38 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_36 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_37 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_43 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_44 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_64 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_63 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_61 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_62 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_68 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_41 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_42 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_69 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_70 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_71 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_72 ;
    wire \FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_73 ;
    wire \FSM_TEST_inst_RAPIDA.N_256_g ;
    wire RST_N_c;
    wire RST_N_c_i;
    wire divisor_inst_counter_0;
    wire clk_continuous_fast;
    wire divisor_inst_counter_1;
    wire \FSM_TEST_inst_RAPIDA.N_100_li ;
    wire \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIKIU51Z0Z_1 ;
    wire \FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z2 ;
    wire \FSM_TEST_inst_RAPIDA.N_123_0 ;
    wire clk_out_RNI3LEM;
    wire \FSM_TEST_inst_RAPIDA.current_stateZ0Z_0 ;
    wire \FSM_TEST_inst_RAPIDA.current_stateZ0Z_1 ;
    wire clk_pll_1;
    wire RST_N_c_i_g;
    wire \config_register_latched_dec_inst.STATCNF_0 ;
    wire STATCNF_i_0;
    wire _gnd_net_;

    defparam \top_pll_inst.top_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \top_pll_inst.top_pll_inst .TEST_MODE=1'b0;
    defparam \top_pll_inst.top_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \top_pll_inst.top_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \top_pll_inst.top_pll_inst .FILTER_RANGE=3'b001;
    defparam \top_pll_inst.top_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \top_pll_inst.top_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \top_pll_inst.top_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \top_pll_inst.top_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \top_pll_inst.top_pll_inst .DIVR=4'b0000;
    defparam \top_pll_inst.top_pll_inst .DIVQ=3'b110;
    defparam \top_pll_inst.top_pll_inst .DIVF=7'b0111111;
    defparam \top_pll_inst.top_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \top_pll_inst.top_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__4904),
            .RESETB(N__12104),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_pll_1));
    IO_PAD CLK_ibuf_iopad (
            .OE(N__12279),
            .DIN(N__12278),
            .DOUT(N__12277),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_preio (
            .PADOEN(N__12279),
            .PADOUT(N__12278),
            .PADIN(N__12277),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD xor_out_stat_obuf_iopad (
            .OE(N__12270),
            .DIN(N__12269),
            .DOUT(N__12268),
            .PACKAGEPIN(xor_out_stat));
    defparam xor_out_stat_obuf_preio.NEG_TRIGGER=1'b0;
    defparam xor_out_stat_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO xor_out_stat_obuf_preio (
            .PADOEN(N__12270),
            .PADOUT(N__12269),
            .PADIN(N__12268),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10442),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_output_obuf_iopad (
            .OE(N__12261),
            .DIN(N__12260),
            .DOUT(N__12259),
            .PACKAGEPIN(clk_output));
    defparam clk_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO clk_output_obuf_preio (
            .PADOEN(N__12261),
            .PADOUT(N__12260),
            .PADIN(N__12259),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8303),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s13_obuf_iopad (
            .OE(N__12252),
            .DIN(N__12251),
            .DOUT(N__12250),
            .PACKAGEPIN(s13));
    defparam s13_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s13_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s13_obuf_preio (
            .PADOEN(N__12252),
            .PADOUT(N__12251),
            .PADIN(N__12250),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6812),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sel_output_obuf_iopad (
            .OE(N__12243),
            .DIN(N__12242),
            .DOUT(N__12241),
            .PACKAGEPIN(sel_output));
    defparam sel_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sel_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sel_output_obuf_preio (
            .PADOEN(N__12243),
            .PADOUT(N__12242),
            .PADIN(N__12241),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10112),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD xor_out_dyn_obuf_iopad (
            .OE(N__12234),
            .DIN(N__12233),
            .DOUT(N__12232),
            .PACKAGEPIN(xor_out_dyn));
    defparam xor_out_dyn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam xor_out_dyn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO xor_out_dyn_obuf_preio (
            .PADOEN(N__12234),
            .PADOUT(N__12233),
            .PADIN(N__12232),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4958),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s12_obuf_iopad (
            .OE(N__12225),
            .DIN(N__12224),
            .DOUT(N__12223),
            .PACKAGEPIN(s12));
    defparam s12_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s12_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s12_obuf_preio (
            .PADOEN(N__12225),
            .PADOUT(N__12224),
            .PADIN(N__12223),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6854),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD miso_input_ibuf_iopad (
            .OE(N__12216),
            .DIN(N__12215),
            .DOUT(N__12214),
            .PACKAGEPIN(miso_input));
    defparam miso_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam miso_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO miso_input_ibuf_preio (
            .PADOEN(N__12216),
            .PADOUT(N__12215),
            .PADIN(N__12214),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(miso_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RST_N_ibuf_iopad (
            .OE(N__12207),
            .DIN(N__12206),
            .DOUT(N__12205),
            .PACKAGEPIN(RST_N));
    defparam RST_N_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RST_N_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RST_N_ibuf_preio (
            .PADOEN(N__12207),
            .PADOUT(N__12206),
            .PADIN(N__12205),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RST_N_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD mosi_output_obuf_iopad (
            .OE(N__12198),
            .DIN(N__12197),
            .DOUT(N__12196),
            .PACKAGEPIN(mosi_output));
    defparam mosi_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam mosi_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO mosi_output_obuf_preio (
            .PADOEN(N__12198),
            .PADOUT(N__12197),
            .PADIN(N__12196),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8027),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s14_obuf_iopad (
            .OE(N__12189),
            .DIN(N__12188),
            .DOUT(N__12187),
            .PACKAGEPIN(s14));
    defparam s14_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s14_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s14_obuf_preio (
            .PADOEN(N__12189),
            .PADOUT(N__12188),
            .PADIN(N__12187),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7985),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2841 (
            .O(N__12170),
            .I(N__12167));
    LocalMux I__2840 (
            .O(N__12167),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_71 ));
    InMux I__2839 (
            .O(N__12164),
            .I(N__12161));
    LocalMux I__2838 (
            .O(N__12161),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_72 ));
    InMux I__2837 (
            .O(N__12158),
            .I(N__12155));
    LocalMux I__2836 (
            .O(N__12155),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_73 ));
    CEMux I__2835 (
            .O(N__12152),
            .I(N__12110));
    CEMux I__2834 (
            .O(N__12151),
            .I(N__12110));
    CEMux I__2833 (
            .O(N__12150),
            .I(N__12110));
    CEMux I__2832 (
            .O(N__12149),
            .I(N__12110));
    CEMux I__2831 (
            .O(N__12148),
            .I(N__12110));
    CEMux I__2830 (
            .O(N__12147),
            .I(N__12110));
    CEMux I__2829 (
            .O(N__12146),
            .I(N__12110));
    CEMux I__2828 (
            .O(N__12145),
            .I(N__12110));
    CEMux I__2827 (
            .O(N__12144),
            .I(N__12110));
    CEMux I__2826 (
            .O(N__12143),
            .I(N__12110));
    CEMux I__2825 (
            .O(N__12142),
            .I(N__12110));
    CEMux I__2824 (
            .O(N__12141),
            .I(N__12110));
    CEMux I__2823 (
            .O(N__12140),
            .I(N__12110));
    CEMux I__2822 (
            .O(N__12139),
            .I(N__12110));
    GlobalMux I__2821 (
            .O(N__12110),
            .I(N__12107));
    gio2CtrlBuf I__2820 (
            .O(N__12107),
            .I(\FSM_TEST_inst_RAPIDA.N_256_g ));
    IoInMux I__2819 (
            .O(N__12104),
            .I(N__12101));
    LocalMux I__2818 (
            .O(N__12101),
            .I(N__12098));
    IoSpan4Mux I__2817 (
            .O(N__12098),
            .I(N__12092));
    InMux I__2816 (
            .O(N__12097),
            .I(N__12089));
    InMux I__2815 (
            .O(N__12096),
            .I(N__12084));
    InMux I__2814 (
            .O(N__12095),
            .I(N__12084));
    Span4Mux_s3_v I__2813 (
            .O(N__12092),
            .I(N__12078));
    LocalMux I__2812 (
            .O(N__12089),
            .I(N__12075));
    LocalMux I__2811 (
            .O(N__12084),
            .I(N__12072));
    CascadeMux I__2810 (
            .O(N__12083),
            .I(N__12067));
    CascadeMux I__2809 (
            .O(N__12082),
            .I(N__12064));
    CascadeMux I__2808 (
            .O(N__12081),
            .I(N__12059));
    Sp12to4 I__2807 (
            .O(N__12078),
            .I(N__12056));
    Span4Mux_v I__2806 (
            .O(N__12075),
            .I(N__12053));
    Span4Mux_v I__2805 (
            .O(N__12072),
            .I(N__12050));
    InMux I__2804 (
            .O(N__12071),
            .I(N__12035));
    InMux I__2803 (
            .O(N__12070),
            .I(N__12035));
    InMux I__2802 (
            .O(N__12067),
            .I(N__12035));
    InMux I__2801 (
            .O(N__12064),
            .I(N__12035));
    InMux I__2800 (
            .O(N__12063),
            .I(N__12035));
    InMux I__2799 (
            .O(N__12062),
            .I(N__12035));
    InMux I__2798 (
            .O(N__12059),
            .I(N__12035));
    Span12Mux_v I__2797 (
            .O(N__12056),
            .I(N__12025));
    Sp12to4 I__2796 (
            .O(N__12053),
            .I(N__12025));
    Sp12to4 I__2795 (
            .O(N__12050),
            .I(N__12025));
    LocalMux I__2794 (
            .O(N__12035),
            .I(N__12025));
    InMux I__2793 (
            .O(N__12034),
            .I(N__12022));
    Span12Mux_h I__2792 (
            .O(N__12025),
            .I(N__12019));
    LocalMux I__2791 (
            .O(N__12022),
            .I(N__12016));
    Span12Mux_v I__2790 (
            .O(N__12019),
            .I(N__12011));
    Span12Mux_h I__2789 (
            .O(N__12016),
            .I(N__12011));
    Odrv12 I__2788 (
            .O(N__12011),
            .I(RST_N_c));
    IoInMux I__2787 (
            .O(N__12008),
            .I(N__12005));
    LocalMux I__2786 (
            .O(N__12005),
            .I(N__12002));
    Odrv12 I__2785 (
            .O(N__12002),
            .I(RST_N_c_i));
    InMux I__2784 (
            .O(N__11999),
            .I(N__11993));
    InMux I__2783 (
            .O(N__11998),
            .I(N__11985));
    InMux I__2782 (
            .O(N__11997),
            .I(N__11985));
    InMux I__2781 (
            .O(N__11996),
            .I(N__11985));
    LocalMux I__2780 (
            .O(N__11993),
            .I(N__11982));
    InMux I__2779 (
            .O(N__11992),
            .I(N__11979));
    LocalMux I__2778 (
            .O(N__11985),
            .I(divisor_inst_counter_0));
    Odrv4 I__2777 (
            .O(N__11982),
            .I(divisor_inst_counter_0));
    LocalMux I__2776 (
            .O(N__11979),
            .I(divisor_inst_counter_0));
    InMux I__2775 (
            .O(N__11972),
            .I(N__11969));
    LocalMux I__2774 (
            .O(N__11969),
            .I(N__11965));
    InMux I__2773 (
            .O(N__11968),
            .I(N__11961));
    Span4Mux_v I__2772 (
            .O(N__11965),
            .I(N__11957));
    InMux I__2771 (
            .O(N__11964),
            .I(N__11954));
    LocalMux I__2770 (
            .O(N__11961),
            .I(N__11951));
    InMux I__2769 (
            .O(N__11960),
            .I(N__11948));
    Odrv4 I__2768 (
            .O(N__11957),
            .I(clk_continuous_fast));
    LocalMux I__2767 (
            .O(N__11954),
            .I(clk_continuous_fast));
    Odrv4 I__2766 (
            .O(N__11951),
            .I(clk_continuous_fast));
    LocalMux I__2765 (
            .O(N__11948),
            .I(clk_continuous_fast));
    CascadeMux I__2764 (
            .O(N__11939),
            .I(N__11936));
    InMux I__2763 (
            .O(N__11936),
            .I(N__11931));
    InMux I__2762 (
            .O(N__11935),
            .I(N__11925));
    InMux I__2761 (
            .O(N__11934),
            .I(N__11925));
    LocalMux I__2760 (
            .O(N__11931),
            .I(N__11922));
    InMux I__2759 (
            .O(N__11930),
            .I(N__11919));
    LocalMux I__2758 (
            .O(N__11925),
            .I(divisor_inst_counter_1));
    Odrv4 I__2757 (
            .O(N__11922),
            .I(divisor_inst_counter_1));
    LocalMux I__2756 (
            .O(N__11919),
            .I(divisor_inst_counter_1));
    InMux I__2755 (
            .O(N__11912),
            .I(N__11905));
    InMux I__2754 (
            .O(N__11911),
            .I(N__11902));
    InMux I__2753 (
            .O(N__11910),
            .I(N__11895));
    InMux I__2752 (
            .O(N__11909),
            .I(N__11895));
    InMux I__2751 (
            .O(N__11908),
            .I(N__11895));
    LocalMux I__2750 (
            .O(N__11905),
            .I(N__11892));
    LocalMux I__2749 (
            .O(N__11902),
            .I(\FSM_TEST_inst_RAPIDA.N_100_li ));
    LocalMux I__2748 (
            .O(N__11895),
            .I(\FSM_TEST_inst_RAPIDA.N_100_li ));
    Odrv12 I__2747 (
            .O(N__11892),
            .I(\FSM_TEST_inst_RAPIDA.N_100_li ));
    IoInMux I__2746 (
            .O(N__11885),
            .I(N__11882));
    LocalMux I__2745 (
            .O(N__11882),
            .I(N__11879));
    Span12Mux_s5_v I__2744 (
            .O(N__11879),
            .I(N__11876));
    Odrv12 I__2743 (
            .O(N__11876),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIKIU51Z0Z_1 ));
    InMux I__2742 (
            .O(N__11873),
            .I(N__11854));
    InMux I__2741 (
            .O(N__11872),
            .I(N__11854));
    InMux I__2740 (
            .O(N__11871),
            .I(N__11854));
    CascadeMux I__2739 (
            .O(N__11870),
            .I(N__11848));
    InMux I__2738 (
            .O(N__11869),
            .I(N__11836));
    InMux I__2737 (
            .O(N__11868),
            .I(N__11836));
    InMux I__2736 (
            .O(N__11867),
            .I(N__11836));
    InMux I__2735 (
            .O(N__11866),
            .I(N__11836));
    InMux I__2734 (
            .O(N__11865),
            .I(N__11836));
    InMux I__2733 (
            .O(N__11864),
            .I(N__11821));
    InMux I__2732 (
            .O(N__11863),
            .I(N__11818));
    InMux I__2731 (
            .O(N__11862),
            .I(N__11813));
    InMux I__2730 (
            .O(N__11861),
            .I(N__11813));
    LocalMux I__2729 (
            .O(N__11854),
            .I(N__11807));
    InMux I__2728 (
            .O(N__11853),
            .I(N__11802));
    InMux I__2727 (
            .O(N__11852),
            .I(N__11802));
    InMux I__2726 (
            .O(N__11851),
            .I(N__11795));
    InMux I__2725 (
            .O(N__11848),
            .I(N__11795));
    InMux I__2724 (
            .O(N__11847),
            .I(N__11795));
    LocalMux I__2723 (
            .O(N__11836),
            .I(N__11792));
    InMux I__2722 (
            .O(N__11835),
            .I(N__11781));
    InMux I__2721 (
            .O(N__11834),
            .I(N__11781));
    InMux I__2720 (
            .O(N__11833),
            .I(N__11781));
    InMux I__2719 (
            .O(N__11832),
            .I(N__11781));
    InMux I__2718 (
            .O(N__11831),
            .I(N__11781));
    InMux I__2717 (
            .O(N__11830),
            .I(N__11772));
    InMux I__2716 (
            .O(N__11829),
            .I(N__11772));
    InMux I__2715 (
            .O(N__11828),
            .I(N__11772));
    InMux I__2714 (
            .O(N__11827),
            .I(N__11772));
    InMux I__2713 (
            .O(N__11826),
            .I(N__11765));
    InMux I__2712 (
            .O(N__11825),
            .I(N__11765));
    InMux I__2711 (
            .O(N__11824),
            .I(N__11765));
    LocalMux I__2710 (
            .O(N__11821),
            .I(N__11760));
    LocalMux I__2709 (
            .O(N__11818),
            .I(N__11760));
    LocalMux I__2708 (
            .O(N__11813),
            .I(N__11757));
    InMux I__2707 (
            .O(N__11812),
            .I(N__11750));
    InMux I__2706 (
            .O(N__11811),
            .I(N__11750));
    InMux I__2705 (
            .O(N__11810),
            .I(N__11750));
    Span4Mux_h I__2704 (
            .O(N__11807),
            .I(N__11744));
    LocalMux I__2703 (
            .O(N__11802),
            .I(N__11744));
    LocalMux I__2702 (
            .O(N__11795),
            .I(N__11741));
    Span4Mux_v I__2701 (
            .O(N__11792),
            .I(N__11736));
    LocalMux I__2700 (
            .O(N__11781),
            .I(N__11736));
    LocalMux I__2699 (
            .O(N__11772),
            .I(N__11731));
    LocalMux I__2698 (
            .O(N__11765),
            .I(N__11731));
    Span4Mux_v I__2697 (
            .O(N__11760),
            .I(N__11724));
    Span4Mux_h I__2696 (
            .O(N__11757),
            .I(N__11724));
    LocalMux I__2695 (
            .O(N__11750),
            .I(N__11724));
    CascadeMux I__2694 (
            .O(N__11749),
            .I(N__11720));
    Span4Mux_v I__2693 (
            .O(N__11744),
            .I(N__11717));
    Span4Mux_h I__2692 (
            .O(N__11741),
            .I(N__11712));
    Span4Mux_h I__2691 (
            .O(N__11736),
            .I(N__11712));
    Span4Mux_v I__2690 (
            .O(N__11731),
            .I(N__11707));
    Span4Mux_h I__2689 (
            .O(N__11724),
            .I(N__11707));
    InMux I__2688 (
            .O(N__11723),
            .I(N__11704));
    InMux I__2687 (
            .O(N__11720),
            .I(N__11701));
    Odrv4 I__2686 (
            .O(N__11717),
            .I(\FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z2 ));
    Odrv4 I__2685 (
            .O(N__11712),
            .I(\FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z2 ));
    Odrv4 I__2684 (
            .O(N__11707),
            .I(\FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z2 ));
    LocalMux I__2683 (
            .O(N__11704),
            .I(\FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z2 ));
    LocalMux I__2682 (
            .O(N__11701),
            .I(\FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z2 ));
    CascadeMux I__2681 (
            .O(N__11690),
            .I(N__11686));
    InMux I__2680 (
            .O(N__11689),
            .I(N__11675));
    InMux I__2679 (
            .O(N__11686),
            .I(N__11675));
    InMux I__2678 (
            .O(N__11685),
            .I(N__11675));
    InMux I__2677 (
            .O(N__11684),
            .I(N__11675));
    LocalMux I__2676 (
            .O(N__11675),
            .I(N__11672));
    Span4Mux_h I__2675 (
            .O(N__11672),
            .I(N__11667));
    InMux I__2674 (
            .O(N__11671),
            .I(N__11662));
    InMux I__2673 (
            .O(N__11670),
            .I(N__11662));
    Odrv4 I__2672 (
            .O(N__11667),
            .I(\FSM_TEST_inst_RAPIDA.N_123_0 ));
    LocalMux I__2671 (
            .O(N__11662),
            .I(\FSM_TEST_inst_RAPIDA.N_123_0 ));
    CascadeMux I__2670 (
            .O(N__11657),
            .I(N__11652));
    InMux I__2669 (
            .O(N__11656),
            .I(N__11646));
    InMux I__2668 (
            .O(N__11655),
            .I(N__11643));
    InMux I__2667 (
            .O(N__11652),
            .I(N__11639));
    InMux I__2666 (
            .O(N__11651),
            .I(N__11636));
    InMux I__2665 (
            .O(N__11650),
            .I(N__11633));
    InMux I__2664 (
            .O(N__11649),
            .I(N__11630));
    LocalMux I__2663 (
            .O(N__11646),
            .I(N__11625));
    LocalMux I__2662 (
            .O(N__11643),
            .I(N__11625));
    CEMux I__2661 (
            .O(N__11642),
            .I(N__11610));
    LocalMux I__2660 (
            .O(N__11639),
            .I(N__11603));
    LocalMux I__2659 (
            .O(N__11636),
            .I(N__11603));
    LocalMux I__2658 (
            .O(N__11633),
            .I(N__11603));
    LocalMux I__2657 (
            .O(N__11630),
            .I(N__11600));
    Span4Mux_h I__2656 (
            .O(N__11625),
            .I(N__11595));
    InMux I__2655 (
            .O(N__11624),
            .I(N__11584));
    InMux I__2654 (
            .O(N__11623),
            .I(N__11584));
    InMux I__2653 (
            .O(N__11622),
            .I(N__11584));
    InMux I__2652 (
            .O(N__11621),
            .I(N__11584));
    InMux I__2651 (
            .O(N__11620),
            .I(N__11584));
    InMux I__2650 (
            .O(N__11619),
            .I(N__11581));
    InMux I__2649 (
            .O(N__11618),
            .I(N__11578));
    InMux I__2648 (
            .O(N__11617),
            .I(N__11567));
    InMux I__2647 (
            .O(N__11616),
            .I(N__11567));
    InMux I__2646 (
            .O(N__11615),
            .I(N__11567));
    InMux I__2645 (
            .O(N__11614),
            .I(N__11567));
    InMux I__2644 (
            .O(N__11613),
            .I(N__11567));
    LocalMux I__2643 (
            .O(N__11610),
            .I(N__11562));
    Span4Mux_v I__2642 (
            .O(N__11603),
            .I(N__11562));
    Span4Mux_h I__2641 (
            .O(N__11600),
            .I(N__11559));
    InMux I__2640 (
            .O(N__11599),
            .I(N__11556));
    InMux I__2639 (
            .O(N__11598),
            .I(N__11553));
    Odrv4 I__2638 (
            .O(N__11595),
            .I(clk_out_RNI3LEM));
    LocalMux I__2637 (
            .O(N__11584),
            .I(clk_out_RNI3LEM));
    LocalMux I__2636 (
            .O(N__11581),
            .I(clk_out_RNI3LEM));
    LocalMux I__2635 (
            .O(N__11578),
            .I(clk_out_RNI3LEM));
    LocalMux I__2634 (
            .O(N__11567),
            .I(clk_out_RNI3LEM));
    Odrv4 I__2633 (
            .O(N__11562),
            .I(clk_out_RNI3LEM));
    Odrv4 I__2632 (
            .O(N__11559),
            .I(clk_out_RNI3LEM));
    LocalMux I__2631 (
            .O(N__11556),
            .I(clk_out_RNI3LEM));
    LocalMux I__2630 (
            .O(N__11553),
            .I(clk_out_RNI3LEM));
    InMux I__2629 (
            .O(N__11534),
            .I(N__11490));
    InMux I__2628 (
            .O(N__11533),
            .I(N__11439));
    InMux I__2627 (
            .O(N__11532),
            .I(N__11439));
    InMux I__2626 (
            .O(N__11531),
            .I(N__11439));
    InMux I__2625 (
            .O(N__11530),
            .I(N__11439));
    InMux I__2624 (
            .O(N__11529),
            .I(N__11439));
    InMux I__2623 (
            .O(N__11528),
            .I(N__11439));
    InMux I__2622 (
            .O(N__11527),
            .I(N__11439));
    InMux I__2621 (
            .O(N__11526),
            .I(N__11426));
    InMux I__2620 (
            .O(N__11525),
            .I(N__11426));
    InMux I__2619 (
            .O(N__11524),
            .I(N__11426));
    InMux I__2618 (
            .O(N__11523),
            .I(N__11426));
    InMux I__2617 (
            .O(N__11522),
            .I(N__11426));
    InMux I__2616 (
            .O(N__11521),
            .I(N__11426));
    InMux I__2615 (
            .O(N__11520),
            .I(N__11409));
    InMux I__2614 (
            .O(N__11519),
            .I(N__11409));
    InMux I__2613 (
            .O(N__11518),
            .I(N__11409));
    InMux I__2612 (
            .O(N__11517),
            .I(N__11409));
    InMux I__2611 (
            .O(N__11516),
            .I(N__11409));
    InMux I__2610 (
            .O(N__11515),
            .I(N__11409));
    InMux I__2609 (
            .O(N__11514),
            .I(N__11409));
    InMux I__2608 (
            .O(N__11513),
            .I(N__11409));
    InMux I__2607 (
            .O(N__11512),
            .I(N__11402));
    InMux I__2606 (
            .O(N__11511),
            .I(N__11402));
    InMux I__2605 (
            .O(N__11510),
            .I(N__11402));
    InMux I__2604 (
            .O(N__11509),
            .I(N__11385));
    InMux I__2603 (
            .O(N__11508),
            .I(N__11385));
    InMux I__2602 (
            .O(N__11507),
            .I(N__11385));
    InMux I__2601 (
            .O(N__11506),
            .I(N__11385));
    InMux I__2600 (
            .O(N__11505),
            .I(N__11385));
    InMux I__2599 (
            .O(N__11504),
            .I(N__11385));
    InMux I__2598 (
            .O(N__11503),
            .I(N__11385));
    InMux I__2597 (
            .O(N__11502),
            .I(N__11385));
    InMux I__2596 (
            .O(N__11501),
            .I(N__11370));
    InMux I__2595 (
            .O(N__11500),
            .I(N__11370));
    InMux I__2594 (
            .O(N__11499),
            .I(N__11370));
    InMux I__2593 (
            .O(N__11498),
            .I(N__11370));
    InMux I__2592 (
            .O(N__11497),
            .I(N__11370));
    InMux I__2591 (
            .O(N__11496),
            .I(N__11370));
    InMux I__2590 (
            .O(N__11495),
            .I(N__11370));
    InMux I__2589 (
            .O(N__11494),
            .I(N__11361));
    InMux I__2588 (
            .O(N__11493),
            .I(N__11361));
    LocalMux I__2587 (
            .O(N__11490),
            .I(N__11358));
    InMux I__2586 (
            .O(N__11489),
            .I(N__11343));
    InMux I__2585 (
            .O(N__11488),
            .I(N__11343));
    InMux I__2584 (
            .O(N__11487),
            .I(N__11343));
    InMux I__2583 (
            .O(N__11486),
            .I(N__11343));
    InMux I__2582 (
            .O(N__11485),
            .I(N__11343));
    InMux I__2581 (
            .O(N__11484),
            .I(N__11343));
    InMux I__2580 (
            .O(N__11483),
            .I(N__11343));
    InMux I__2579 (
            .O(N__11482),
            .I(N__11330));
    InMux I__2578 (
            .O(N__11481),
            .I(N__11330));
    InMux I__2577 (
            .O(N__11480),
            .I(N__11330));
    InMux I__2576 (
            .O(N__11479),
            .I(N__11330));
    InMux I__2575 (
            .O(N__11478),
            .I(N__11330));
    InMux I__2574 (
            .O(N__11477),
            .I(N__11330));
    InMux I__2573 (
            .O(N__11476),
            .I(N__11323));
    InMux I__2572 (
            .O(N__11475),
            .I(N__11323));
    InMux I__2571 (
            .O(N__11474),
            .I(N__11323));
    InMux I__2570 (
            .O(N__11473),
            .I(N__11308));
    InMux I__2569 (
            .O(N__11472),
            .I(N__11308));
    InMux I__2568 (
            .O(N__11471),
            .I(N__11308));
    InMux I__2567 (
            .O(N__11470),
            .I(N__11308));
    InMux I__2566 (
            .O(N__11469),
            .I(N__11308));
    InMux I__2565 (
            .O(N__11468),
            .I(N__11308));
    InMux I__2564 (
            .O(N__11467),
            .I(N__11308));
    InMux I__2563 (
            .O(N__11466),
            .I(N__11305));
    InMux I__2562 (
            .O(N__11465),
            .I(N__11296));
    InMux I__2561 (
            .O(N__11464),
            .I(N__11296));
    InMux I__2560 (
            .O(N__11463),
            .I(N__11296));
    InMux I__2559 (
            .O(N__11462),
            .I(N__11296));
    InMux I__2558 (
            .O(N__11461),
            .I(N__11291));
    InMux I__2557 (
            .O(N__11460),
            .I(N__11291));
    InMux I__2556 (
            .O(N__11459),
            .I(N__11288));
    InMux I__2555 (
            .O(N__11458),
            .I(N__11243));
    InMux I__2554 (
            .O(N__11457),
            .I(N__11243));
    InMux I__2553 (
            .O(N__11456),
            .I(N__11243));
    InMux I__2552 (
            .O(N__11455),
            .I(N__11243));
    InMux I__2551 (
            .O(N__11454),
            .I(N__11243));
    LocalMux I__2550 (
            .O(N__11439),
            .I(N__11230));
    LocalMux I__2549 (
            .O(N__11426),
            .I(N__11230));
    LocalMux I__2548 (
            .O(N__11409),
            .I(N__11230));
    LocalMux I__2547 (
            .O(N__11402),
            .I(N__11230));
    LocalMux I__2546 (
            .O(N__11385),
            .I(N__11230));
    LocalMux I__2545 (
            .O(N__11370),
            .I(N__11230));
    InMux I__2544 (
            .O(N__11369),
            .I(N__11221));
    InMux I__2543 (
            .O(N__11368),
            .I(N__11221));
    InMux I__2542 (
            .O(N__11367),
            .I(N__11221));
    InMux I__2541 (
            .O(N__11366),
            .I(N__11221));
    LocalMux I__2540 (
            .O(N__11361),
            .I(N__11214));
    Span4Mux_v I__2539 (
            .O(N__11358),
            .I(N__11214));
    LocalMux I__2538 (
            .O(N__11343),
            .I(N__11199));
    LocalMux I__2537 (
            .O(N__11330),
            .I(N__11199));
    LocalMux I__2536 (
            .O(N__11323),
            .I(N__11199));
    LocalMux I__2535 (
            .O(N__11308),
            .I(N__11199));
    LocalMux I__2534 (
            .O(N__11305),
            .I(N__11199));
    LocalMux I__2533 (
            .O(N__11296),
            .I(N__11199));
    LocalMux I__2532 (
            .O(N__11291),
            .I(N__11199));
    LocalMux I__2531 (
            .O(N__11288),
            .I(N__11196));
    InMux I__2530 (
            .O(N__11287),
            .I(N__11188));
    InMux I__2529 (
            .O(N__11286),
            .I(N__11188));
    InMux I__2528 (
            .O(N__11285),
            .I(N__11173));
    InMux I__2527 (
            .O(N__11284),
            .I(N__11173));
    InMux I__2526 (
            .O(N__11283),
            .I(N__11173));
    InMux I__2525 (
            .O(N__11282),
            .I(N__11173));
    InMux I__2524 (
            .O(N__11281),
            .I(N__11173));
    InMux I__2523 (
            .O(N__11280),
            .I(N__11173));
    InMux I__2522 (
            .O(N__11279),
            .I(N__11173));
    InMux I__2521 (
            .O(N__11278),
            .I(N__11158));
    InMux I__2520 (
            .O(N__11277),
            .I(N__11158));
    InMux I__2519 (
            .O(N__11276),
            .I(N__11158));
    InMux I__2518 (
            .O(N__11275),
            .I(N__11158));
    InMux I__2517 (
            .O(N__11274),
            .I(N__11158));
    InMux I__2516 (
            .O(N__11273),
            .I(N__11158));
    InMux I__2515 (
            .O(N__11272),
            .I(N__11158));
    InMux I__2514 (
            .O(N__11271),
            .I(N__11153));
    InMux I__2513 (
            .O(N__11270),
            .I(N__11153));
    InMux I__2512 (
            .O(N__11269),
            .I(N__11150));
    InMux I__2511 (
            .O(N__11268),
            .I(N__11140));
    InMux I__2510 (
            .O(N__11267),
            .I(N__11140));
    InMux I__2509 (
            .O(N__11266),
            .I(N__11140));
    InMux I__2508 (
            .O(N__11265),
            .I(N__11125));
    InMux I__2507 (
            .O(N__11264),
            .I(N__11125));
    InMux I__2506 (
            .O(N__11263),
            .I(N__11125));
    InMux I__2505 (
            .O(N__11262),
            .I(N__11125));
    InMux I__2504 (
            .O(N__11261),
            .I(N__11125));
    InMux I__2503 (
            .O(N__11260),
            .I(N__11125));
    InMux I__2502 (
            .O(N__11259),
            .I(N__11125));
    InMux I__2501 (
            .O(N__11258),
            .I(N__11114));
    InMux I__2500 (
            .O(N__11257),
            .I(N__11114));
    InMux I__2499 (
            .O(N__11256),
            .I(N__11114));
    InMux I__2498 (
            .O(N__11255),
            .I(N__11114));
    InMux I__2497 (
            .O(N__11254),
            .I(N__11114));
    LocalMux I__2496 (
            .O(N__11243),
            .I(N__11107));
    Span4Mux_v I__2495 (
            .O(N__11230),
            .I(N__11107));
    LocalMux I__2494 (
            .O(N__11221),
            .I(N__11107));
    InMux I__2493 (
            .O(N__11220),
            .I(N__11104));
    InMux I__2492 (
            .O(N__11219),
            .I(N__11101));
    Span4Mux_h I__2491 (
            .O(N__11214),
            .I(N__11094));
    Span4Mux_v I__2490 (
            .O(N__11199),
            .I(N__11094));
    Span4Mux_v I__2489 (
            .O(N__11196),
            .I(N__11094));
    InMux I__2488 (
            .O(N__11195),
            .I(N__11087));
    InMux I__2487 (
            .O(N__11194),
            .I(N__11087));
    InMux I__2486 (
            .O(N__11193),
            .I(N__11087));
    LocalMux I__2485 (
            .O(N__11188),
            .I(N__11078));
    LocalMux I__2484 (
            .O(N__11173),
            .I(N__11078));
    LocalMux I__2483 (
            .O(N__11158),
            .I(N__11078));
    LocalMux I__2482 (
            .O(N__11153),
            .I(N__11078));
    LocalMux I__2481 (
            .O(N__11150),
            .I(N__11075));
    InMux I__2480 (
            .O(N__11149),
            .I(N__11068));
    InMux I__2479 (
            .O(N__11148),
            .I(N__11068));
    InMux I__2478 (
            .O(N__11147),
            .I(N__11068));
    LocalMux I__2477 (
            .O(N__11140),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_0 ));
    LocalMux I__2476 (
            .O(N__11125),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_0 ));
    LocalMux I__2475 (
            .O(N__11114),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_0 ));
    Odrv4 I__2474 (
            .O(N__11107),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_0 ));
    LocalMux I__2473 (
            .O(N__11104),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_0 ));
    LocalMux I__2472 (
            .O(N__11101),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_0 ));
    Odrv4 I__2471 (
            .O(N__11094),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_0 ));
    LocalMux I__2470 (
            .O(N__11087),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_0 ));
    Odrv4 I__2469 (
            .O(N__11078),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_0 ));
    Odrv4 I__2468 (
            .O(N__11075),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_0 ));
    LocalMux I__2467 (
            .O(N__11068),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_0 ));
    InMux I__2466 (
            .O(N__11045),
            .I(N__11034));
    InMux I__2465 (
            .O(N__11044),
            .I(N__11034));
    InMux I__2464 (
            .O(N__11043),
            .I(N__11011));
    InMux I__2463 (
            .O(N__11042),
            .I(N__11011));
    InMux I__2462 (
            .O(N__11041),
            .I(N__11011));
    InMux I__2461 (
            .O(N__11040),
            .I(N__11011));
    InMux I__2460 (
            .O(N__11039),
            .I(N__11011));
    LocalMux I__2459 (
            .O(N__11034),
            .I(N__11008));
    InMux I__2458 (
            .O(N__11033),
            .I(N__11005));
    InMux I__2457 (
            .O(N__11032),
            .I(N__10996));
    InMux I__2456 (
            .O(N__11031),
            .I(N__10989));
    InMux I__2455 (
            .O(N__11030),
            .I(N__10989));
    InMux I__2454 (
            .O(N__11029),
            .I(N__10989));
    InMux I__2453 (
            .O(N__11028),
            .I(N__10982));
    InMux I__2452 (
            .O(N__11027),
            .I(N__10982));
    InMux I__2451 (
            .O(N__11026),
            .I(N__10982));
    InMux I__2450 (
            .O(N__11025),
            .I(N__10973));
    InMux I__2449 (
            .O(N__11024),
            .I(N__10973));
    InMux I__2448 (
            .O(N__11023),
            .I(N__10973));
    InMux I__2447 (
            .O(N__11022),
            .I(N__10973));
    LocalMux I__2446 (
            .O(N__11011),
            .I(N__10964));
    Span4Mux_h I__2445 (
            .O(N__11008),
            .I(N__10959));
    LocalMux I__2444 (
            .O(N__11005),
            .I(N__10959));
    InMux I__2443 (
            .O(N__11004),
            .I(N__10952));
    InMux I__2442 (
            .O(N__11003),
            .I(N__10952));
    InMux I__2441 (
            .O(N__11002),
            .I(N__10952));
    InMux I__2440 (
            .O(N__11001),
            .I(N__10945));
    InMux I__2439 (
            .O(N__11000),
            .I(N__10945));
    InMux I__2438 (
            .O(N__10999),
            .I(N__10945));
    LocalMux I__2437 (
            .O(N__10996),
            .I(N__10934));
    LocalMux I__2436 (
            .O(N__10989),
            .I(N__10934));
    LocalMux I__2435 (
            .O(N__10982),
            .I(N__10934));
    LocalMux I__2434 (
            .O(N__10973),
            .I(N__10934));
    InMux I__2433 (
            .O(N__10972),
            .I(N__10923));
    InMux I__2432 (
            .O(N__10971),
            .I(N__10923));
    InMux I__2431 (
            .O(N__10970),
            .I(N__10923));
    InMux I__2430 (
            .O(N__10969),
            .I(N__10923));
    InMux I__2429 (
            .O(N__10968),
            .I(N__10923));
    CascadeMux I__2428 (
            .O(N__10967),
            .I(N__10920));
    Span4Mux_h I__2427 (
            .O(N__10964),
            .I(N__10911));
    Span4Mux_h I__2426 (
            .O(N__10959),
            .I(N__10911));
    LocalMux I__2425 (
            .O(N__10952),
            .I(N__10911));
    LocalMux I__2424 (
            .O(N__10945),
            .I(N__10911));
    InMux I__2423 (
            .O(N__10944),
            .I(N__10906));
    InMux I__2422 (
            .O(N__10943),
            .I(N__10906));
    Span4Mux_v I__2421 (
            .O(N__10934),
            .I(N__10901));
    LocalMux I__2420 (
            .O(N__10923),
            .I(N__10901));
    InMux I__2419 (
            .O(N__10920),
            .I(N__10898));
    Odrv4 I__2418 (
            .O(N__10911),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_1 ));
    LocalMux I__2417 (
            .O(N__10906),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_1 ));
    Odrv4 I__2416 (
            .O(N__10901),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_1 ));
    LocalMux I__2415 (
            .O(N__10898),
            .I(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_1 ));
    ClkMux I__2414 (
            .O(N__10889),
            .I(N__10676));
    ClkMux I__2413 (
            .O(N__10888),
            .I(N__10676));
    ClkMux I__2412 (
            .O(N__10887),
            .I(N__10676));
    ClkMux I__2411 (
            .O(N__10886),
            .I(N__10676));
    ClkMux I__2410 (
            .O(N__10885),
            .I(N__10676));
    ClkMux I__2409 (
            .O(N__10884),
            .I(N__10676));
    ClkMux I__2408 (
            .O(N__10883),
            .I(N__10676));
    ClkMux I__2407 (
            .O(N__10882),
            .I(N__10676));
    ClkMux I__2406 (
            .O(N__10881),
            .I(N__10676));
    ClkMux I__2405 (
            .O(N__10880),
            .I(N__10676));
    ClkMux I__2404 (
            .O(N__10879),
            .I(N__10676));
    ClkMux I__2403 (
            .O(N__10878),
            .I(N__10676));
    ClkMux I__2402 (
            .O(N__10877),
            .I(N__10676));
    ClkMux I__2401 (
            .O(N__10876),
            .I(N__10676));
    ClkMux I__2400 (
            .O(N__10875),
            .I(N__10676));
    ClkMux I__2399 (
            .O(N__10874),
            .I(N__10676));
    ClkMux I__2398 (
            .O(N__10873),
            .I(N__10676));
    ClkMux I__2397 (
            .O(N__10872),
            .I(N__10676));
    ClkMux I__2396 (
            .O(N__10871),
            .I(N__10676));
    ClkMux I__2395 (
            .O(N__10870),
            .I(N__10676));
    ClkMux I__2394 (
            .O(N__10869),
            .I(N__10676));
    ClkMux I__2393 (
            .O(N__10868),
            .I(N__10676));
    ClkMux I__2392 (
            .O(N__10867),
            .I(N__10676));
    ClkMux I__2391 (
            .O(N__10866),
            .I(N__10676));
    ClkMux I__2390 (
            .O(N__10865),
            .I(N__10676));
    ClkMux I__2389 (
            .O(N__10864),
            .I(N__10676));
    ClkMux I__2388 (
            .O(N__10863),
            .I(N__10676));
    ClkMux I__2387 (
            .O(N__10862),
            .I(N__10676));
    ClkMux I__2386 (
            .O(N__10861),
            .I(N__10676));
    ClkMux I__2385 (
            .O(N__10860),
            .I(N__10676));
    ClkMux I__2384 (
            .O(N__10859),
            .I(N__10676));
    ClkMux I__2383 (
            .O(N__10858),
            .I(N__10676));
    ClkMux I__2382 (
            .O(N__10857),
            .I(N__10676));
    ClkMux I__2381 (
            .O(N__10856),
            .I(N__10676));
    ClkMux I__2380 (
            .O(N__10855),
            .I(N__10676));
    ClkMux I__2379 (
            .O(N__10854),
            .I(N__10676));
    ClkMux I__2378 (
            .O(N__10853),
            .I(N__10676));
    ClkMux I__2377 (
            .O(N__10852),
            .I(N__10676));
    ClkMux I__2376 (
            .O(N__10851),
            .I(N__10676));
    ClkMux I__2375 (
            .O(N__10850),
            .I(N__10676));
    ClkMux I__2374 (
            .O(N__10849),
            .I(N__10676));
    ClkMux I__2373 (
            .O(N__10848),
            .I(N__10676));
    ClkMux I__2372 (
            .O(N__10847),
            .I(N__10676));
    ClkMux I__2371 (
            .O(N__10846),
            .I(N__10676));
    ClkMux I__2370 (
            .O(N__10845),
            .I(N__10676));
    ClkMux I__2369 (
            .O(N__10844),
            .I(N__10676));
    ClkMux I__2368 (
            .O(N__10843),
            .I(N__10676));
    ClkMux I__2367 (
            .O(N__10842),
            .I(N__10676));
    ClkMux I__2366 (
            .O(N__10841),
            .I(N__10676));
    ClkMux I__2365 (
            .O(N__10840),
            .I(N__10676));
    ClkMux I__2364 (
            .O(N__10839),
            .I(N__10676));
    ClkMux I__2363 (
            .O(N__10838),
            .I(N__10676));
    ClkMux I__2362 (
            .O(N__10837),
            .I(N__10676));
    ClkMux I__2361 (
            .O(N__10836),
            .I(N__10676));
    ClkMux I__2360 (
            .O(N__10835),
            .I(N__10676));
    ClkMux I__2359 (
            .O(N__10834),
            .I(N__10676));
    ClkMux I__2358 (
            .O(N__10833),
            .I(N__10676));
    ClkMux I__2357 (
            .O(N__10832),
            .I(N__10676));
    ClkMux I__2356 (
            .O(N__10831),
            .I(N__10676));
    ClkMux I__2355 (
            .O(N__10830),
            .I(N__10676));
    ClkMux I__2354 (
            .O(N__10829),
            .I(N__10676));
    ClkMux I__2353 (
            .O(N__10828),
            .I(N__10676));
    ClkMux I__2352 (
            .O(N__10827),
            .I(N__10676));
    ClkMux I__2351 (
            .O(N__10826),
            .I(N__10676));
    ClkMux I__2350 (
            .O(N__10825),
            .I(N__10676));
    ClkMux I__2349 (
            .O(N__10824),
            .I(N__10676));
    ClkMux I__2348 (
            .O(N__10823),
            .I(N__10676));
    ClkMux I__2347 (
            .O(N__10822),
            .I(N__10676));
    ClkMux I__2346 (
            .O(N__10821),
            .I(N__10676));
    ClkMux I__2345 (
            .O(N__10820),
            .I(N__10676));
    ClkMux I__2344 (
            .O(N__10819),
            .I(N__10676));
    GlobalMux I__2343 (
            .O(N__10676),
            .I(clk_pll_1));
    SRMux I__2342 (
            .O(N__10673),
            .I(N__10460));
    SRMux I__2341 (
            .O(N__10672),
            .I(N__10460));
    SRMux I__2340 (
            .O(N__10671),
            .I(N__10460));
    SRMux I__2339 (
            .O(N__10670),
            .I(N__10460));
    SRMux I__2338 (
            .O(N__10669),
            .I(N__10460));
    SRMux I__2337 (
            .O(N__10668),
            .I(N__10460));
    SRMux I__2336 (
            .O(N__10667),
            .I(N__10460));
    SRMux I__2335 (
            .O(N__10666),
            .I(N__10460));
    SRMux I__2334 (
            .O(N__10665),
            .I(N__10460));
    SRMux I__2333 (
            .O(N__10664),
            .I(N__10460));
    SRMux I__2332 (
            .O(N__10663),
            .I(N__10460));
    SRMux I__2331 (
            .O(N__10662),
            .I(N__10460));
    SRMux I__2330 (
            .O(N__10661),
            .I(N__10460));
    SRMux I__2329 (
            .O(N__10660),
            .I(N__10460));
    SRMux I__2328 (
            .O(N__10659),
            .I(N__10460));
    SRMux I__2327 (
            .O(N__10658),
            .I(N__10460));
    SRMux I__2326 (
            .O(N__10657),
            .I(N__10460));
    SRMux I__2325 (
            .O(N__10656),
            .I(N__10460));
    SRMux I__2324 (
            .O(N__10655),
            .I(N__10460));
    SRMux I__2323 (
            .O(N__10654),
            .I(N__10460));
    SRMux I__2322 (
            .O(N__10653),
            .I(N__10460));
    SRMux I__2321 (
            .O(N__10652),
            .I(N__10460));
    SRMux I__2320 (
            .O(N__10651),
            .I(N__10460));
    SRMux I__2319 (
            .O(N__10650),
            .I(N__10460));
    SRMux I__2318 (
            .O(N__10649),
            .I(N__10460));
    SRMux I__2317 (
            .O(N__10648),
            .I(N__10460));
    SRMux I__2316 (
            .O(N__10647),
            .I(N__10460));
    SRMux I__2315 (
            .O(N__10646),
            .I(N__10460));
    SRMux I__2314 (
            .O(N__10645),
            .I(N__10460));
    SRMux I__2313 (
            .O(N__10644),
            .I(N__10460));
    SRMux I__2312 (
            .O(N__10643),
            .I(N__10460));
    SRMux I__2311 (
            .O(N__10642),
            .I(N__10460));
    SRMux I__2310 (
            .O(N__10641),
            .I(N__10460));
    SRMux I__2309 (
            .O(N__10640),
            .I(N__10460));
    SRMux I__2308 (
            .O(N__10639),
            .I(N__10460));
    SRMux I__2307 (
            .O(N__10638),
            .I(N__10460));
    SRMux I__2306 (
            .O(N__10637),
            .I(N__10460));
    SRMux I__2305 (
            .O(N__10636),
            .I(N__10460));
    SRMux I__2304 (
            .O(N__10635),
            .I(N__10460));
    SRMux I__2303 (
            .O(N__10634),
            .I(N__10460));
    SRMux I__2302 (
            .O(N__10633),
            .I(N__10460));
    SRMux I__2301 (
            .O(N__10632),
            .I(N__10460));
    SRMux I__2300 (
            .O(N__10631),
            .I(N__10460));
    SRMux I__2299 (
            .O(N__10630),
            .I(N__10460));
    SRMux I__2298 (
            .O(N__10629),
            .I(N__10460));
    SRMux I__2297 (
            .O(N__10628),
            .I(N__10460));
    SRMux I__2296 (
            .O(N__10627),
            .I(N__10460));
    SRMux I__2295 (
            .O(N__10626),
            .I(N__10460));
    SRMux I__2294 (
            .O(N__10625),
            .I(N__10460));
    SRMux I__2293 (
            .O(N__10624),
            .I(N__10460));
    SRMux I__2292 (
            .O(N__10623),
            .I(N__10460));
    SRMux I__2291 (
            .O(N__10622),
            .I(N__10460));
    SRMux I__2290 (
            .O(N__10621),
            .I(N__10460));
    SRMux I__2289 (
            .O(N__10620),
            .I(N__10460));
    SRMux I__2288 (
            .O(N__10619),
            .I(N__10460));
    SRMux I__2287 (
            .O(N__10618),
            .I(N__10460));
    SRMux I__2286 (
            .O(N__10617),
            .I(N__10460));
    SRMux I__2285 (
            .O(N__10616),
            .I(N__10460));
    SRMux I__2284 (
            .O(N__10615),
            .I(N__10460));
    SRMux I__2283 (
            .O(N__10614),
            .I(N__10460));
    SRMux I__2282 (
            .O(N__10613),
            .I(N__10460));
    SRMux I__2281 (
            .O(N__10612),
            .I(N__10460));
    SRMux I__2280 (
            .O(N__10611),
            .I(N__10460));
    SRMux I__2279 (
            .O(N__10610),
            .I(N__10460));
    SRMux I__2278 (
            .O(N__10609),
            .I(N__10460));
    SRMux I__2277 (
            .O(N__10608),
            .I(N__10460));
    SRMux I__2276 (
            .O(N__10607),
            .I(N__10460));
    SRMux I__2275 (
            .O(N__10606),
            .I(N__10460));
    SRMux I__2274 (
            .O(N__10605),
            .I(N__10460));
    SRMux I__2273 (
            .O(N__10604),
            .I(N__10460));
    SRMux I__2272 (
            .O(N__10603),
            .I(N__10460));
    GlobalMux I__2271 (
            .O(N__10460),
            .I(N__10457));
    gio2CtrlBuf I__2270 (
            .O(N__10457),
            .I(RST_N_c_i_g));
    InMux I__2269 (
            .O(N__10454),
            .I(N__10451));
    LocalMux I__2268 (
            .O(N__10451),
            .I(N__10448));
    Span4Mux_h I__2267 (
            .O(N__10448),
            .I(N__10445));
    Odrv4 I__2266 (
            .O(N__10445),
            .I(\config_register_latched_dec_inst.STATCNF_0 ));
    IoInMux I__2265 (
            .O(N__10442),
            .I(N__10439));
    LocalMux I__2264 (
            .O(N__10439),
            .I(N__10436));
    Span4Mux_s3_h I__2263 (
            .O(N__10436),
            .I(N__10433));
    Span4Mux_h I__2262 (
            .O(N__10433),
            .I(N__10430));
    Span4Mux_h I__2261 (
            .O(N__10430),
            .I(N__10427));
    Odrv4 I__2260 (
            .O(N__10427),
            .I(STATCNF_i_0));
    InMux I__2259 (
            .O(N__10424),
            .I(N__10421));
    LocalMux I__2258 (
            .O(N__10421),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_37 ));
    InMux I__2257 (
            .O(N__10418),
            .I(N__10415));
    LocalMux I__2256 (
            .O(N__10415),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_43 ));
    InMux I__2255 (
            .O(N__10412),
            .I(N__10409));
    LocalMux I__2254 (
            .O(N__10409),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_44 ));
    InMux I__2253 (
            .O(N__10406),
            .I(N__10403));
    LocalMux I__2252 (
            .O(N__10403),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_64 ));
    InMux I__2251 (
            .O(N__10400),
            .I(N__10397));
    LocalMux I__2250 (
            .O(N__10397),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_63 ));
    InMux I__2249 (
            .O(N__10394),
            .I(N__10391));
    LocalMux I__2248 (
            .O(N__10391),
            .I(N__10388));
    Odrv4 I__2247 (
            .O(N__10388),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_61 ));
    InMux I__2246 (
            .O(N__10385),
            .I(N__10382));
    LocalMux I__2245 (
            .O(N__10382),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_62 ));
    InMux I__2244 (
            .O(N__10379),
            .I(N__10376));
    LocalMux I__2243 (
            .O(N__10376),
            .I(N__10373));
    Odrv4 I__2242 (
            .O(N__10373),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_68 ));
    InMux I__2241 (
            .O(N__10370),
            .I(N__10367));
    LocalMux I__2240 (
            .O(N__10367),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_41 ));
    CascadeMux I__2239 (
            .O(N__10364),
            .I(N__10361));
    InMux I__2238 (
            .O(N__10361),
            .I(N__10358));
    LocalMux I__2237 (
            .O(N__10358),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_42 ));
    InMux I__2236 (
            .O(N__10355),
            .I(N__10352));
    LocalMux I__2235 (
            .O(N__10352),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_69 ));
    InMux I__2234 (
            .O(N__10349),
            .I(N__10346));
    LocalMux I__2233 (
            .O(N__10346),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_70 ));
    CascadeMux I__2232 (
            .O(N__10343),
            .I(N__10321));
    CascadeMux I__2231 (
            .O(N__10342),
            .I(N__10318));
    CascadeMux I__2230 (
            .O(N__10341),
            .I(N__10315));
    InMux I__2229 (
            .O(N__10340),
            .I(N__10291));
    InMux I__2228 (
            .O(N__10339),
            .I(N__10291));
    InMux I__2227 (
            .O(N__10338),
            .I(N__10291));
    InMux I__2226 (
            .O(N__10337),
            .I(N__10291));
    InMux I__2225 (
            .O(N__10336),
            .I(N__10291));
    InMux I__2224 (
            .O(N__10335),
            .I(N__10291));
    InMux I__2223 (
            .O(N__10334),
            .I(N__10291));
    InMux I__2222 (
            .O(N__10333),
            .I(N__10282));
    InMux I__2221 (
            .O(N__10332),
            .I(N__10282));
    InMux I__2220 (
            .O(N__10331),
            .I(N__10282));
    InMux I__2219 (
            .O(N__10330),
            .I(N__10282));
    InMux I__2218 (
            .O(N__10329),
            .I(N__10279));
    InMux I__2217 (
            .O(N__10328),
            .I(N__10272));
    InMux I__2216 (
            .O(N__10327),
            .I(N__10272));
    InMux I__2215 (
            .O(N__10326),
            .I(N__10272));
    InMux I__2214 (
            .O(N__10325),
            .I(N__10267));
    InMux I__2213 (
            .O(N__10324),
            .I(N__10267));
    InMux I__2212 (
            .O(N__10321),
            .I(N__10260));
    InMux I__2211 (
            .O(N__10318),
            .I(N__10260));
    InMux I__2210 (
            .O(N__10315),
            .I(N__10260));
    CascadeMux I__2209 (
            .O(N__10314),
            .I(N__10255));
    CascadeMux I__2208 (
            .O(N__10313),
            .I(N__10252));
    CascadeMux I__2207 (
            .O(N__10312),
            .I(N__10249));
    CascadeMux I__2206 (
            .O(N__10311),
            .I(N__10246));
    InMux I__2205 (
            .O(N__10310),
            .I(N__10232));
    InMux I__2204 (
            .O(N__10309),
            .I(N__10232));
    InMux I__2203 (
            .O(N__10308),
            .I(N__10232));
    InMux I__2202 (
            .O(N__10307),
            .I(N__10232));
    InMux I__2201 (
            .O(N__10306),
            .I(N__10232));
    LocalMux I__2200 (
            .O(N__10291),
            .I(N__10227));
    LocalMux I__2199 (
            .O(N__10282),
            .I(N__10227));
    LocalMux I__2198 (
            .O(N__10279),
            .I(N__10218));
    LocalMux I__2197 (
            .O(N__10272),
            .I(N__10218));
    LocalMux I__2196 (
            .O(N__10267),
            .I(N__10218));
    LocalMux I__2195 (
            .O(N__10260),
            .I(N__10218));
    InMux I__2194 (
            .O(N__10259),
            .I(N__10215));
    InMux I__2193 (
            .O(N__10258),
            .I(N__10202));
    InMux I__2192 (
            .O(N__10255),
            .I(N__10202));
    InMux I__2191 (
            .O(N__10252),
            .I(N__10202));
    InMux I__2190 (
            .O(N__10249),
            .I(N__10202));
    InMux I__2189 (
            .O(N__10246),
            .I(N__10202));
    InMux I__2188 (
            .O(N__10245),
            .I(N__10202));
    InMux I__2187 (
            .O(N__10244),
            .I(N__10199));
    CascadeMux I__2186 (
            .O(N__10243),
            .I(N__10196));
    LocalMux I__2185 (
            .O(N__10232),
            .I(N__10193));
    Span4Mux_v I__2184 (
            .O(N__10227),
            .I(N__10188));
    Span4Mux_v I__2183 (
            .O(N__10218),
            .I(N__10188));
    LocalMux I__2182 (
            .O(N__10215),
            .I(N__10181));
    LocalMux I__2181 (
            .O(N__10202),
            .I(N__10181));
    LocalMux I__2180 (
            .O(N__10199),
            .I(N__10181));
    InMux I__2179 (
            .O(N__10196),
            .I(N__10178));
    Odrv4 I__2178 (
            .O(N__10193),
            .I(\FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z1 ));
    Odrv4 I__2177 (
            .O(N__10188),
            .I(\FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z1 ));
    Odrv4 I__2176 (
            .O(N__10181),
            .I(\FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z1 ));
    LocalMux I__2175 (
            .O(N__10178),
            .I(\FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z1 ));
    InMux I__2174 (
            .O(N__10169),
            .I(N__10166));
    LocalMux I__2173 (
            .O(N__10166),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_11 ));
    InMux I__2172 (
            .O(N__10163),
            .I(N__10160));
    LocalMux I__2171 (
            .O(N__10160),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_12 ));
    InMux I__2170 (
            .O(N__10157),
            .I(N__10154));
    LocalMux I__2169 (
            .O(N__10154),
            .I(N__10150));
    CascadeMux I__2168 (
            .O(N__10153),
            .I(N__10146));
    Span4Mux_v I__2167 (
            .O(N__10150),
            .I(N__10143));
    InMux I__2166 (
            .O(N__10149),
            .I(N__10140));
    InMux I__2165 (
            .O(N__10146),
            .I(N__10137));
    Odrv4 I__2164 (
            .O(N__10143),
            .I(\config_register_latched_dec_inst.STATSRZ0Z_0 ));
    LocalMux I__2163 (
            .O(N__10140),
            .I(\config_register_latched_dec_inst.STATSRZ0Z_0 ));
    LocalMux I__2162 (
            .O(N__10137),
            .I(\config_register_latched_dec_inst.STATSRZ0Z_0 ));
    CascadeMux I__2161 (
            .O(N__10130),
            .I(N__10127));
    InMux I__2160 (
            .O(N__10127),
            .I(N__10124));
    LocalMux I__2159 (
            .O(N__10124),
            .I(N__10120));
    InMux I__2158 (
            .O(N__10123),
            .I(N__10117));
    Odrv4 I__2157 (
            .O(N__10120),
            .I(\config_register_latched_dec_inst.STATCNF_1Z0Z_0 ));
    LocalMux I__2156 (
            .O(N__10117),
            .I(\config_register_latched_dec_inst.STATCNF_1Z0Z_0 ));
    IoInMux I__2155 (
            .O(N__10112),
            .I(N__10109));
    LocalMux I__2154 (
            .O(N__10109),
            .I(N__10106));
    IoSpan4Mux I__2153 (
            .O(N__10106),
            .I(N__10102));
    CascadeMux I__2152 (
            .O(N__10105),
            .I(N__10099));
    Span4Mux_s2_h I__2151 (
            .O(N__10102),
            .I(N__10095));
    InMux I__2150 (
            .O(N__10099),
            .I(N__10089));
    InMux I__2149 (
            .O(N__10098),
            .I(N__10089));
    Span4Mux_h I__2148 (
            .O(N__10095),
            .I(N__10075));
    InMux I__2147 (
            .O(N__10094),
            .I(N__10064));
    LocalMux I__2146 (
            .O(N__10089),
            .I(N__10061));
    InMux I__2145 (
            .O(N__10088),
            .I(N__10050));
    InMux I__2144 (
            .O(N__10087),
            .I(N__10050));
    InMux I__2143 (
            .O(N__10086),
            .I(N__10050));
    InMux I__2142 (
            .O(N__10085),
            .I(N__10050));
    InMux I__2141 (
            .O(N__10084),
            .I(N__10050));
    InMux I__2140 (
            .O(N__10083),
            .I(N__10047));
    InMux I__2139 (
            .O(N__10082),
            .I(N__10042));
    InMux I__2138 (
            .O(N__10081),
            .I(N__10042));
    InMux I__2137 (
            .O(N__10080),
            .I(N__10035));
    InMux I__2136 (
            .O(N__10079),
            .I(N__10035));
    InMux I__2135 (
            .O(N__10078),
            .I(N__10035));
    Sp12to4 I__2134 (
            .O(N__10075),
            .I(N__10032));
    InMux I__2133 (
            .O(N__10074),
            .I(N__10021));
    InMux I__2132 (
            .O(N__10073),
            .I(N__10021));
    InMux I__2131 (
            .O(N__10072),
            .I(N__10021));
    InMux I__2130 (
            .O(N__10071),
            .I(N__10021));
    InMux I__2129 (
            .O(N__10070),
            .I(N__10021));
    InMux I__2128 (
            .O(N__10069),
            .I(N__10014));
    InMux I__2127 (
            .O(N__10068),
            .I(N__10014));
    InMux I__2126 (
            .O(N__10067),
            .I(N__10014));
    LocalMux I__2125 (
            .O(N__10064),
            .I(N__10011));
    Span4Mux_v I__2124 (
            .O(N__10061),
            .I(N__10008));
    LocalMux I__2123 (
            .O(N__10050),
            .I(N__9999));
    LocalMux I__2122 (
            .O(N__10047),
            .I(N__9999));
    LocalMux I__2121 (
            .O(N__10042),
            .I(N__9999));
    LocalMux I__2120 (
            .O(N__10035),
            .I(N__9999));
    Span12Mux_h I__2119 (
            .O(N__10032),
            .I(N__9996));
    LocalMux I__2118 (
            .O(N__10021),
            .I(N__9991));
    LocalMux I__2117 (
            .O(N__10014),
            .I(N__9991));
    Span4Mux_v I__2116 (
            .O(N__10011),
            .I(N__9984));
    Span4Mux_h I__2115 (
            .O(N__10008),
            .I(N__9984));
    Span4Mux_v I__2114 (
            .O(N__9999),
            .I(N__9984));
    Odrv12 I__2113 (
            .O(N__9996),
            .I(sel_output_c));
    Odrv12 I__2112 (
            .O(N__9991),
            .I(sel_output_c));
    Odrv4 I__2111 (
            .O(N__9984),
            .I(sel_output_c));
    CascadeMux I__2110 (
            .O(N__9977),
            .I(N__9974));
    InMux I__2109 (
            .O(N__9974),
            .I(N__9967));
    InMux I__2108 (
            .O(N__9973),
            .I(N__9964));
    InMux I__2107 (
            .O(N__9972),
            .I(N__9961));
    InMux I__2106 (
            .O(N__9971),
            .I(N__9956));
    InMux I__2105 (
            .O(N__9970),
            .I(N__9956));
    LocalMux I__2104 (
            .O(N__9967),
            .I(N__9951));
    LocalMux I__2103 (
            .O(N__9964),
            .I(N__9951));
    LocalMux I__2102 (
            .O(N__9961),
            .I(N__9948));
    LocalMux I__2101 (
            .O(N__9956),
            .I(\FSM_TEST_inst_RAPIDA.counter_dinZ0Z_2 ));
    Odrv4 I__2100 (
            .O(N__9951),
            .I(\FSM_TEST_inst_RAPIDA.counter_dinZ0Z_2 ));
    Odrv12 I__2099 (
            .O(N__9948),
            .I(\FSM_TEST_inst_RAPIDA.counter_dinZ0Z_2 ));
    InMux I__2098 (
            .O(N__9941),
            .I(N__9937));
    CascadeMux I__2097 (
            .O(N__9940),
            .I(N__9933));
    LocalMux I__2096 (
            .O(N__9937),
            .I(N__9928));
    InMux I__2095 (
            .O(N__9936),
            .I(N__9925));
    InMux I__2094 (
            .O(N__9933),
            .I(N__9918));
    InMux I__2093 (
            .O(N__9932),
            .I(N__9918));
    InMux I__2092 (
            .O(N__9931),
            .I(N__9918));
    Odrv12 I__2091 (
            .O(N__9928),
            .I(\FSM_TEST_inst_RAPIDA.counter_dinZ1Z_1 ));
    LocalMux I__2090 (
            .O(N__9925),
            .I(\FSM_TEST_inst_RAPIDA.counter_dinZ1Z_1 ));
    LocalMux I__2089 (
            .O(N__9918),
            .I(\FSM_TEST_inst_RAPIDA.counter_dinZ1Z_1 ));
    CascadeMux I__2088 (
            .O(N__9911),
            .I(N__9906));
    CascadeMux I__2087 (
            .O(N__9910),
            .I(N__9903));
    CascadeMux I__2086 (
            .O(N__9909),
            .I(N__9900));
    InMux I__2085 (
            .O(N__9906),
            .I(N__9897));
    InMux I__2084 (
            .O(N__9903),
            .I(N__9894));
    InMux I__2083 (
            .O(N__9900),
            .I(N__9891));
    LocalMux I__2082 (
            .O(N__9897),
            .I(N__9888));
    LocalMux I__2081 (
            .O(N__9894),
            .I(\FSM_TEST_inst_RAPIDA.counter_dinZ0Z_3 ));
    LocalMux I__2080 (
            .O(N__9891),
            .I(\FSM_TEST_inst_RAPIDA.counter_dinZ0Z_3 ));
    Odrv12 I__2079 (
            .O(N__9888),
            .I(\FSM_TEST_inst_RAPIDA.counter_dinZ0Z_3 ));
    InMux I__2078 (
            .O(N__9881),
            .I(N__9874));
    InMux I__2077 (
            .O(N__9880),
            .I(N__9866));
    InMux I__2076 (
            .O(N__9879),
            .I(N__9866));
    InMux I__2075 (
            .O(N__9878),
            .I(N__9866));
    InMux I__2074 (
            .O(N__9877),
            .I(N__9863));
    LocalMux I__2073 (
            .O(N__9874),
            .I(N__9860));
    InMux I__2072 (
            .O(N__9873),
            .I(N__9857));
    LocalMux I__2071 (
            .O(N__9866),
            .I(N__9854));
    LocalMux I__2070 (
            .O(N__9863),
            .I(\FSM_TEST_inst_RAPIDA.counter_dinZ0Z_0 ));
    Odrv4 I__2069 (
            .O(N__9860),
            .I(\FSM_TEST_inst_RAPIDA.counter_dinZ0Z_0 ));
    LocalMux I__2068 (
            .O(N__9857),
            .I(\FSM_TEST_inst_RAPIDA.counter_dinZ0Z_0 ));
    Odrv4 I__2067 (
            .O(N__9854),
            .I(\FSM_TEST_inst_RAPIDA.counter_dinZ0Z_0 ));
    InMux I__2066 (
            .O(N__9845),
            .I(N__9842));
    LocalMux I__2065 (
            .O(N__9842),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_66 ));
    InMux I__2064 (
            .O(N__9839),
            .I(N__9836));
    LocalMux I__2063 (
            .O(N__9836),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_67 ));
    InMux I__2062 (
            .O(N__9833),
            .I(N__9830));
    LocalMux I__2061 (
            .O(N__9830),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_45 ));
    InMux I__2060 (
            .O(N__9827),
            .I(N__9824));
    LocalMux I__2059 (
            .O(N__9824),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_38 ));
    InMux I__2058 (
            .O(N__9821),
            .I(N__9818));
    LocalMux I__2057 (
            .O(N__9818),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_36 ));
    InMux I__2056 (
            .O(N__9815),
            .I(N__9812));
    LocalMux I__2055 (
            .O(N__9812),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_48 ));
    InMux I__2054 (
            .O(N__9809),
            .I(N__9806));
    LocalMux I__2053 (
            .O(N__9806),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_49 ));
    InMux I__2052 (
            .O(N__9803),
            .I(N__9800));
    LocalMux I__2051 (
            .O(N__9800),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_33 ));
    InMux I__2050 (
            .O(N__9797),
            .I(N__9794));
    LocalMux I__2049 (
            .O(N__9794),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_34 ));
    InMux I__2048 (
            .O(N__9791),
            .I(N__9788));
    LocalMux I__2047 (
            .O(N__9788),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_10 ));
    InMux I__2046 (
            .O(N__9785),
            .I(N__9782));
    LocalMux I__2045 (
            .O(N__9782),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_74 ));
    InMux I__2044 (
            .O(N__9779),
            .I(N__9776));
    LocalMux I__2043 (
            .O(N__9776),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_13 ));
    InMux I__2042 (
            .O(N__9773),
            .I(N__9770));
    LocalMux I__2041 (
            .O(N__9770),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_14 ));
    InMux I__2040 (
            .O(N__9767),
            .I(N__9764));
    LocalMux I__2039 (
            .O(N__9764),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_15 ));
    InMux I__2038 (
            .O(N__9761),
            .I(N__9758));
    LocalMux I__2037 (
            .O(N__9758),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_16 ));
    InMux I__2036 (
            .O(N__9755),
            .I(N__9752));
    LocalMux I__2035 (
            .O(N__9752),
            .I(N__9749));
    Odrv4 I__2034 (
            .O(N__9749),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_17 ));
    InMux I__2033 (
            .O(N__9746),
            .I(N__9743));
    LocalMux I__2032 (
            .O(N__9743),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_65 ));
    InMux I__2031 (
            .O(N__9740),
            .I(N__9737));
    LocalMux I__2030 (
            .O(N__9737),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_35 ));
    InMux I__2029 (
            .O(N__9734),
            .I(N__9731));
    LocalMux I__2028 (
            .O(N__9731),
            .I(N__9728));
    Odrv4 I__2027 (
            .O(N__9728),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_80 ));
    InMux I__2026 (
            .O(N__9725),
            .I(N__9722));
    LocalMux I__2025 (
            .O(N__9722),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_81 ));
    InMux I__2024 (
            .O(N__9719),
            .I(N__9716));
    LocalMux I__2023 (
            .O(N__9716),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_32 ));
    InMux I__2022 (
            .O(N__9713),
            .I(N__9710));
    LocalMux I__2021 (
            .O(N__9710),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_39 ));
    InMux I__2020 (
            .O(N__9707),
            .I(N__9704));
    LocalMux I__2019 (
            .O(N__9704),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_46 ));
    InMux I__2018 (
            .O(N__9701),
            .I(N__9698));
    LocalMux I__2017 (
            .O(N__9698),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_47 ));
    InMux I__2016 (
            .O(N__9695),
            .I(N__9692));
    LocalMux I__2015 (
            .O(N__9692),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_40 ));
    InMux I__2014 (
            .O(N__9689),
            .I(N__9686));
    LocalMux I__2013 (
            .O(N__9686),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_55 ));
    InMux I__2012 (
            .O(N__9683),
            .I(N__9680));
    LocalMux I__2011 (
            .O(N__9680),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_56 ));
    InMux I__2010 (
            .O(N__9677),
            .I(N__9674));
    LocalMux I__2009 (
            .O(N__9674),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_83 ));
    CascadeMux I__2008 (
            .O(N__9671),
            .I(N__9668));
    InMux I__2007 (
            .O(N__9668),
            .I(N__9665));
    LocalMux I__2006 (
            .O(N__9665),
            .I(N__9662));
    Span4Mux_h I__2005 (
            .O(N__9662),
            .I(N__9659));
    Odrv4 I__2004 (
            .O(N__9659),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_87 ));
    InMux I__2003 (
            .O(N__9656),
            .I(N__9653));
    LocalMux I__2002 (
            .O(N__9653),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_84 ));
    InMux I__2001 (
            .O(N__9650),
            .I(N__9647));
    LocalMux I__2000 (
            .O(N__9647),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_85 ));
    InMux I__1999 (
            .O(N__9644),
            .I(N__9641));
    LocalMux I__1998 (
            .O(N__9641),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_86 ));
    InMux I__1997 (
            .O(N__9638),
            .I(N__9635));
    LocalMux I__1996 (
            .O(N__9635),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_82 ));
    InMux I__1995 (
            .O(N__9632),
            .I(N__9629));
    LocalMux I__1994 (
            .O(N__9629),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_29 ));
    InMux I__1993 (
            .O(N__9626),
            .I(N__9623));
    LocalMux I__1992 (
            .O(N__9623),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_30 ));
    InMux I__1991 (
            .O(N__9620),
            .I(N__9617));
    LocalMux I__1990 (
            .O(N__9617),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_75 ));
    InMux I__1989 (
            .O(N__9614),
            .I(N__9611));
    LocalMux I__1988 (
            .O(N__9611),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_60 ));
    InMux I__1987 (
            .O(N__9608),
            .I(N__9605));
    LocalMux I__1986 (
            .O(N__9605),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_58 ));
    InMux I__1985 (
            .O(N__9602),
            .I(N__9599));
    LocalMux I__1984 (
            .O(N__9599),
            .I(N__9596));
    Odrv4 I__1983 (
            .O(N__9596),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_7 ));
    InMux I__1982 (
            .O(N__9593),
            .I(N__9590));
    LocalMux I__1981 (
            .O(N__9590),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_8 ));
    InMux I__1980 (
            .O(N__9587),
            .I(N__9584));
    LocalMux I__1979 (
            .O(N__9584),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_9 ));
    InMux I__1978 (
            .O(N__9581),
            .I(N__9578));
    LocalMux I__1977 (
            .O(N__9578),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_57 ));
    InMux I__1976 (
            .O(N__9575),
            .I(N__9572));
    LocalMux I__1975 (
            .O(N__9572),
            .I(N__9569));
    Span4Mux_h I__1974 (
            .O(N__9569),
            .I(N__9566));
    Odrv4 I__1973 (
            .O(N__9566),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_79 ));
    InMux I__1972 (
            .O(N__9563),
            .I(N__9557));
    InMux I__1971 (
            .O(N__9562),
            .I(N__9557));
    LocalMux I__1970 (
            .O(N__9557),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_7 ));
    InMux I__1969 (
            .O(N__9554),
            .I(N__9548));
    InMux I__1968 (
            .O(N__9553),
            .I(N__9548));
    LocalMux I__1967 (
            .O(N__9548),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_5 ));
    InMux I__1966 (
            .O(N__9545),
            .I(N__9539));
    InMux I__1965 (
            .O(N__9544),
            .I(N__9539));
    LocalMux I__1964 (
            .O(N__9539),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_6 ));
    InMux I__1963 (
            .O(N__9536),
            .I(N__9532));
    InMux I__1962 (
            .O(N__9535),
            .I(N__9529));
    LocalMux I__1961 (
            .O(N__9532),
            .I(N__9522));
    LocalMux I__1960 (
            .O(N__9529),
            .I(N__9522));
    InMux I__1959 (
            .O(N__9528),
            .I(N__9517));
    InMux I__1958 (
            .O(N__9527),
            .I(N__9517));
    Span4Mux_h I__1957 (
            .O(N__9522),
            .I(N__9514));
    LocalMux I__1956 (
            .O(N__9517),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_8 ));
    Odrv4 I__1955 (
            .O(N__9514),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_8 ));
    CascadeMux I__1954 (
            .O(N__9509),
            .I(N__9506));
    InMux I__1953 (
            .O(N__9506),
            .I(N__9500));
    InMux I__1952 (
            .O(N__9505),
            .I(N__9500));
    LocalMux I__1951 (
            .O(N__9500),
            .I(N__9495));
    InMux I__1950 (
            .O(N__9499),
            .I(N__9492));
    InMux I__1949 (
            .O(N__9498),
            .I(N__9489));
    Span4Mux_h I__1948 (
            .O(N__9495),
            .I(N__9486));
    LocalMux I__1947 (
            .O(N__9492),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_9 ));
    LocalMux I__1946 (
            .O(N__9489),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_9 ));
    Odrv4 I__1945 (
            .O(N__9486),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_9 ));
    CEMux I__1944 (
            .O(N__9479),
            .I(N__9475));
    CEMux I__1943 (
            .O(N__9478),
            .I(N__9472));
    LocalMux I__1942 (
            .O(N__9475),
            .I(N__9469));
    LocalMux I__1941 (
            .O(N__9472),
            .I(N__9466));
    Span4Mux_v I__1940 (
            .O(N__9469),
            .I(N__9463));
    Span4Mux_v I__1939 (
            .O(N__9466),
            .I(N__9460));
    Odrv4 I__1938 (
            .O(N__9463),
            .I(flag_output_0_ret_RNI1E8NZ0Z2));
    Odrv4 I__1937 (
            .O(N__9460),
            .I(flag_output_0_ret_RNI1E8NZ0Z2));
    InMux I__1936 (
            .O(N__9455),
            .I(N__9452));
    LocalMux I__1935 (
            .O(N__9452),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_51 ));
    InMux I__1934 (
            .O(N__9449),
            .I(N__9446));
    LocalMux I__1933 (
            .O(N__9446),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_52 ));
    InMux I__1932 (
            .O(N__9443),
            .I(N__9440));
    LocalMux I__1931 (
            .O(N__9440),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_53 ));
    InMux I__1930 (
            .O(N__9437),
            .I(N__9434));
    LocalMux I__1929 (
            .O(N__9434),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_31 ));
    InMux I__1928 (
            .O(N__9431),
            .I(N__9428));
    LocalMux I__1927 (
            .O(N__9428),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_50 ));
    InMux I__1926 (
            .O(N__9425),
            .I(N__9421));
    CascadeMux I__1925 (
            .O(N__9424),
            .I(N__9415));
    LocalMux I__1924 (
            .O(N__9421),
            .I(N__9408));
    InMux I__1923 (
            .O(N__9420),
            .I(N__9405));
    InMux I__1922 (
            .O(N__9419),
            .I(N__9394));
    InMux I__1921 (
            .O(N__9418),
            .I(N__9394));
    InMux I__1920 (
            .O(N__9415),
            .I(N__9394));
    InMux I__1919 (
            .O(N__9414),
            .I(N__9394));
    InMux I__1918 (
            .O(N__9413),
            .I(N__9394));
    InMux I__1917 (
            .O(N__9412),
            .I(N__9391));
    CascadeMux I__1916 (
            .O(N__9411),
            .I(N__9388));
    Span4Mux_h I__1915 (
            .O(N__9408),
            .I(N__9382));
    LocalMux I__1914 (
            .O(N__9405),
            .I(N__9382));
    LocalMux I__1913 (
            .O(N__9394),
            .I(N__9377));
    LocalMux I__1912 (
            .O(N__9391),
            .I(N__9377));
    InMux I__1911 (
            .O(N__9388),
            .I(N__9374));
    InMux I__1910 (
            .O(N__9387),
            .I(N__9371));
    Span4Mux_v I__1909 (
            .O(N__9382),
            .I(N__9368));
    Span4Mux_h I__1908 (
            .O(N__9377),
            .I(N__9365));
    LocalMux I__1907 (
            .O(N__9374),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fastZ0Z_1 ));
    LocalMux I__1906 (
            .O(N__9371),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fastZ0Z_1 ));
    Odrv4 I__1905 (
            .O(N__9368),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fastZ0Z_1 ));
    Odrv4 I__1904 (
            .O(N__9365),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fastZ0Z_1 ));
    InMux I__1903 (
            .O(N__9356),
            .I(N__9353));
    LocalMux I__1902 (
            .O(N__9353),
            .I(N__9350));
    Odrv12 I__1901 (
            .O(N__9350),
            .I(\FSM_TEST_inst_slow.CLK_uC_6kZ0Z_0 ));
    InMux I__1900 (
            .O(N__9347),
            .I(N__9344));
    LocalMux I__1899 (
            .O(N__9344),
            .I(N__9340));
    InMux I__1898 (
            .O(N__9343),
            .I(N__9337));
    Odrv4 I__1897 (
            .O(N__9340),
            .I(CLK_uC_6l_0));
    LocalMux I__1896 (
            .O(N__9337),
            .I(CLK_uC_6l_0));
    InMux I__1895 (
            .O(N__9332),
            .I(N__9326));
    InMux I__1894 (
            .O(N__9331),
            .I(N__9326));
    LocalMux I__1893 (
            .O(N__9326),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_3 ));
    InMux I__1892 (
            .O(N__9323),
            .I(N__9317));
    InMux I__1891 (
            .O(N__9322),
            .I(N__9317));
    LocalMux I__1890 (
            .O(N__9317),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_4 ));
    InMux I__1889 (
            .O(N__9314),
            .I(N__9310));
    InMux I__1888 (
            .O(N__9313),
            .I(N__9307));
    LocalMux I__1887 (
            .O(N__9310),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_1 ));
    LocalMux I__1886 (
            .O(N__9307),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_1 ));
    InMux I__1885 (
            .O(N__9302),
            .I(N__9296));
    InMux I__1884 (
            .O(N__9301),
            .I(N__9296));
    LocalMux I__1883 (
            .O(N__9296),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_2 ));
    InMux I__1882 (
            .O(N__9293),
            .I(N__9284));
    InMux I__1881 (
            .O(N__9292),
            .I(N__9281));
    InMux I__1880 (
            .O(N__9291),
            .I(N__9270));
    InMux I__1879 (
            .O(N__9290),
            .I(N__9270));
    InMux I__1878 (
            .O(N__9289),
            .I(N__9270));
    InMux I__1877 (
            .O(N__9288),
            .I(N__9270));
    InMux I__1876 (
            .O(N__9287),
            .I(N__9270));
    LocalMux I__1875 (
            .O(N__9284),
            .I(N__9265));
    LocalMux I__1874 (
            .O(N__9281),
            .I(N__9265));
    LocalMux I__1873 (
            .O(N__9270),
            .I(\FSM_TEST_inst_slow.current_state_RNI9C3K2Z0Z_1 ));
    Odrv12 I__1872 (
            .O(N__9265),
            .I(\FSM_TEST_inst_slow.current_state_RNI9C3K2Z0Z_1 ));
    CascadeMux I__1871 (
            .O(N__9260),
            .I(N__9256));
    CascadeMux I__1870 (
            .O(N__9259),
            .I(N__9251));
    InMux I__1869 (
            .O(N__9256),
            .I(N__9247));
    CascadeMux I__1868 (
            .O(N__9255),
            .I(N__9244));
    CascadeMux I__1867 (
            .O(N__9254),
            .I(N__9241));
    InMux I__1866 (
            .O(N__9251),
            .I(N__9236));
    InMux I__1865 (
            .O(N__9250),
            .I(N__9233));
    LocalMux I__1864 (
            .O(N__9247),
            .I(N__9230));
    InMux I__1863 (
            .O(N__9244),
            .I(N__9221));
    InMux I__1862 (
            .O(N__9241),
            .I(N__9221));
    InMux I__1861 (
            .O(N__9240),
            .I(N__9221));
    InMux I__1860 (
            .O(N__9239),
            .I(N__9221));
    LocalMux I__1859 (
            .O(N__9236),
            .I(N__9216));
    LocalMux I__1858 (
            .O(N__9233),
            .I(N__9216));
    Span4Mux_h I__1857 (
            .O(N__9230),
            .I(N__9213));
    LocalMux I__1856 (
            .O(N__9221),
            .I(\FSM_TEST_inst_slow.current_state_d_i_2 ));
    Odrv4 I__1855 (
            .O(N__9216),
            .I(\FSM_TEST_inst_slow.current_state_d_i_2 ));
    Odrv4 I__1854 (
            .O(N__9213),
            .I(\FSM_TEST_inst_slow.current_state_d_i_2 ));
    InMux I__1853 (
            .O(N__9206),
            .I(N__9203));
    LocalMux I__1852 (
            .O(N__9203),
            .I(N__9200));
    Odrv4 I__1851 (
            .O(N__9200),
            .I(\FSM_TEST_inst_slow.counter_stat_cry_4_THRU_CO ));
    CascadeMux I__1850 (
            .O(N__9197),
            .I(N__9193));
    InMux I__1849 (
            .O(N__9196),
            .I(N__9189));
    InMux I__1848 (
            .O(N__9193),
            .I(N__9186));
    InMux I__1847 (
            .O(N__9192),
            .I(N__9183));
    LocalMux I__1846 (
            .O(N__9189),
            .I(N__9175));
    LocalMux I__1845 (
            .O(N__9186),
            .I(N__9175));
    LocalMux I__1844 (
            .O(N__9183),
            .I(N__9175));
    InMux I__1843 (
            .O(N__9182),
            .I(N__9172));
    Span4Mux_h I__1842 (
            .O(N__9175),
            .I(N__9169));
    LocalMux I__1841 (
            .O(N__9172),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_5 ));
    Odrv4 I__1840 (
            .O(N__9169),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_5 ));
    InMux I__1839 (
            .O(N__9164),
            .I(N__9153));
    InMux I__1838 (
            .O(N__9163),
            .I(N__9153));
    InMux I__1837 (
            .O(N__9162),
            .I(N__9153));
    InMux I__1836 (
            .O(N__9161),
            .I(N__9148));
    InMux I__1835 (
            .O(N__9160),
            .I(N__9148));
    LocalMux I__1834 (
            .O(N__9153),
            .I(N__9145));
    LocalMux I__1833 (
            .O(N__9148),
            .I(\divisor_inst_2.counterZ0Z_1 ));
    Odrv4 I__1832 (
            .O(N__9145),
            .I(\divisor_inst_2.counterZ0Z_1 ));
    CascadeMux I__1831 (
            .O(N__9140),
            .I(N__9136));
    CascadeMux I__1830 (
            .O(N__9139),
            .I(N__9131));
    InMux I__1829 (
            .O(N__9136),
            .I(N__9122));
    InMux I__1828 (
            .O(N__9135),
            .I(N__9122));
    InMux I__1827 (
            .O(N__9134),
            .I(N__9122));
    InMux I__1826 (
            .O(N__9131),
            .I(N__9115));
    InMux I__1825 (
            .O(N__9130),
            .I(N__9115));
    InMux I__1824 (
            .O(N__9129),
            .I(N__9115));
    LocalMux I__1823 (
            .O(N__9122),
            .I(\divisor_inst_2.counterZ0Z_0 ));
    LocalMux I__1822 (
            .O(N__9115),
            .I(\divisor_inst_2.counterZ0Z_0 ));
    CascadeMux I__1821 (
            .O(N__9110),
            .I(N__9104));
    CascadeMux I__1820 (
            .O(N__9109),
            .I(N__9101));
    InMux I__1819 (
            .O(N__9108),
            .I(N__9098));
    InMux I__1818 (
            .O(N__9107),
            .I(N__9091));
    InMux I__1817 (
            .O(N__9104),
            .I(N__9091));
    InMux I__1816 (
            .O(N__9101),
            .I(N__9091));
    LocalMux I__1815 (
            .O(N__9098),
            .I(\divisor_inst_2.counterZ0Z_2 ));
    LocalMux I__1814 (
            .O(N__9091),
            .I(\divisor_inst_2.counterZ0Z_2 ));
    CascadeMux I__1813 (
            .O(N__9086),
            .I(N__9082));
    CascadeMux I__1812 (
            .O(N__9085),
            .I(N__9078));
    InMux I__1811 (
            .O(N__9082),
            .I(N__9075));
    InMux I__1810 (
            .O(N__9081),
            .I(N__9072));
    InMux I__1809 (
            .O(N__9078),
            .I(N__9069));
    LocalMux I__1808 (
            .O(N__9075),
            .I(\FSM_TEST_inst_RAPIDA.aux_selection_fast_0 ));
    LocalMux I__1807 (
            .O(N__9072),
            .I(\FSM_TEST_inst_RAPIDA.aux_selection_fast_0 ));
    LocalMux I__1806 (
            .O(N__9069),
            .I(\FSM_TEST_inst_RAPIDA.aux_selection_fast_0 ));
    InMux I__1805 (
            .O(N__9062),
            .I(N__9057));
    InMux I__1804 (
            .O(N__9061),
            .I(N__9052));
    InMux I__1803 (
            .O(N__9060),
            .I(N__9052));
    LocalMux I__1802 (
            .O(N__9057),
            .I(N__9038));
    LocalMux I__1801 (
            .O(N__9052),
            .I(N__9035));
    InMux I__1800 (
            .O(N__9051),
            .I(N__9030));
    InMux I__1799 (
            .O(N__9050),
            .I(N__9030));
    InMux I__1798 (
            .O(N__9049),
            .I(N__8995));
    InMux I__1797 (
            .O(N__9048),
            .I(N__8995));
    InMux I__1796 (
            .O(N__9047),
            .I(N__8995));
    InMux I__1795 (
            .O(N__9046),
            .I(N__8992));
    InMux I__1794 (
            .O(N__9045),
            .I(N__8989));
    InMux I__1793 (
            .O(N__9044),
            .I(N__8947));
    InMux I__1792 (
            .O(N__9043),
            .I(N__8942));
    InMux I__1791 (
            .O(N__9042),
            .I(N__8942));
    InMux I__1790 (
            .O(N__9041),
            .I(N__8927));
    Span4Mux_v I__1789 (
            .O(N__9038),
            .I(N__8920));
    Span4Mux_h I__1788 (
            .O(N__9035),
            .I(N__8920));
    LocalMux I__1787 (
            .O(N__9030),
            .I(N__8920));
    InMux I__1786 (
            .O(N__9029),
            .I(N__8909));
    InMux I__1785 (
            .O(N__9028),
            .I(N__8909));
    InMux I__1784 (
            .O(N__9027),
            .I(N__8909));
    InMux I__1783 (
            .O(N__9026),
            .I(N__8909));
    InMux I__1782 (
            .O(N__9025),
            .I(N__8909));
    InMux I__1781 (
            .O(N__9024),
            .I(N__8898));
    InMux I__1780 (
            .O(N__9023),
            .I(N__8898));
    InMux I__1779 (
            .O(N__9022),
            .I(N__8898));
    InMux I__1778 (
            .O(N__9021),
            .I(N__8898));
    InMux I__1777 (
            .O(N__9020),
            .I(N__8898));
    InMux I__1776 (
            .O(N__9019),
            .I(N__8883));
    InMux I__1775 (
            .O(N__9018),
            .I(N__8883));
    InMux I__1774 (
            .O(N__9017),
            .I(N__8883));
    InMux I__1773 (
            .O(N__9016),
            .I(N__8883));
    InMux I__1772 (
            .O(N__9015),
            .I(N__8883));
    InMux I__1771 (
            .O(N__9014),
            .I(N__8883));
    InMux I__1770 (
            .O(N__9013),
            .I(N__8883));
    InMux I__1769 (
            .O(N__9012),
            .I(N__8880));
    InMux I__1768 (
            .O(N__9011),
            .I(N__8863));
    InMux I__1767 (
            .O(N__9010),
            .I(N__8863));
    InMux I__1766 (
            .O(N__9009),
            .I(N__8863));
    InMux I__1765 (
            .O(N__9008),
            .I(N__8863));
    InMux I__1764 (
            .O(N__9007),
            .I(N__8863));
    InMux I__1763 (
            .O(N__9006),
            .I(N__8863));
    InMux I__1762 (
            .O(N__9005),
            .I(N__8863));
    InMux I__1761 (
            .O(N__9004),
            .I(N__8863));
    InMux I__1760 (
            .O(N__9003),
            .I(N__8858));
    InMux I__1759 (
            .O(N__9002),
            .I(N__8858));
    LocalMux I__1758 (
            .O(N__8995),
            .I(N__8851));
    LocalMux I__1757 (
            .O(N__8992),
            .I(N__8848));
    LocalMux I__1756 (
            .O(N__8989),
            .I(N__8845));
    InMux I__1755 (
            .O(N__8988),
            .I(N__8834));
    InMux I__1754 (
            .O(N__8987),
            .I(N__8834));
    InMux I__1753 (
            .O(N__8986),
            .I(N__8834));
    InMux I__1752 (
            .O(N__8985),
            .I(N__8834));
    InMux I__1751 (
            .O(N__8984),
            .I(N__8834));
    InMux I__1750 (
            .O(N__8983),
            .I(N__8827));
    InMux I__1749 (
            .O(N__8982),
            .I(N__8827));
    InMux I__1748 (
            .O(N__8981),
            .I(N__8827));
    InMux I__1747 (
            .O(N__8980),
            .I(N__8824));
    InMux I__1746 (
            .O(N__8979),
            .I(N__8817));
    InMux I__1745 (
            .O(N__8978),
            .I(N__8817));
    InMux I__1744 (
            .O(N__8977),
            .I(N__8817));
    InMux I__1743 (
            .O(N__8976),
            .I(N__8804));
    InMux I__1742 (
            .O(N__8975),
            .I(N__8804));
    InMux I__1741 (
            .O(N__8974),
            .I(N__8804));
    InMux I__1740 (
            .O(N__8973),
            .I(N__8804));
    InMux I__1739 (
            .O(N__8972),
            .I(N__8804));
    InMux I__1738 (
            .O(N__8971),
            .I(N__8804));
    InMux I__1737 (
            .O(N__8970),
            .I(N__8789));
    InMux I__1736 (
            .O(N__8969),
            .I(N__8789));
    InMux I__1735 (
            .O(N__8968),
            .I(N__8789));
    InMux I__1734 (
            .O(N__8967),
            .I(N__8789));
    InMux I__1733 (
            .O(N__8966),
            .I(N__8789));
    InMux I__1732 (
            .O(N__8965),
            .I(N__8789));
    InMux I__1731 (
            .O(N__8964),
            .I(N__8789));
    InMux I__1730 (
            .O(N__8963),
            .I(N__8778));
    InMux I__1729 (
            .O(N__8962),
            .I(N__8778));
    InMux I__1728 (
            .O(N__8961),
            .I(N__8778));
    InMux I__1727 (
            .O(N__8960),
            .I(N__8778));
    InMux I__1726 (
            .O(N__8959),
            .I(N__8778));
    InMux I__1725 (
            .O(N__8958),
            .I(N__8769));
    InMux I__1724 (
            .O(N__8957),
            .I(N__8769));
    InMux I__1723 (
            .O(N__8956),
            .I(N__8769));
    InMux I__1722 (
            .O(N__8955),
            .I(N__8769));
    InMux I__1721 (
            .O(N__8954),
            .I(N__8765));
    InMux I__1720 (
            .O(N__8953),
            .I(N__8756));
    InMux I__1719 (
            .O(N__8952),
            .I(N__8756));
    InMux I__1718 (
            .O(N__8951),
            .I(N__8756));
    InMux I__1717 (
            .O(N__8950),
            .I(N__8756));
    LocalMux I__1716 (
            .O(N__8947),
            .I(N__8751));
    LocalMux I__1715 (
            .O(N__8942),
            .I(N__8751));
    InMux I__1714 (
            .O(N__8941),
            .I(N__8742));
    InMux I__1713 (
            .O(N__8940),
            .I(N__8742));
    InMux I__1712 (
            .O(N__8939),
            .I(N__8742));
    InMux I__1711 (
            .O(N__8938),
            .I(N__8742));
    InMux I__1710 (
            .O(N__8937),
            .I(N__8725));
    InMux I__1709 (
            .O(N__8936),
            .I(N__8725));
    InMux I__1708 (
            .O(N__8935),
            .I(N__8725));
    InMux I__1707 (
            .O(N__8934),
            .I(N__8725));
    InMux I__1706 (
            .O(N__8933),
            .I(N__8725));
    InMux I__1705 (
            .O(N__8932),
            .I(N__8725));
    InMux I__1704 (
            .O(N__8931),
            .I(N__8725));
    InMux I__1703 (
            .O(N__8930),
            .I(N__8725));
    LocalMux I__1702 (
            .O(N__8927),
            .I(N__8698));
    Span4Mux_h I__1701 (
            .O(N__8920),
            .I(N__8698));
    LocalMux I__1700 (
            .O(N__8909),
            .I(N__8698));
    LocalMux I__1699 (
            .O(N__8898),
            .I(N__8698));
    LocalMux I__1698 (
            .O(N__8883),
            .I(N__8698));
    LocalMux I__1697 (
            .O(N__8880),
            .I(N__8695));
    LocalMux I__1696 (
            .O(N__8863),
            .I(N__8690));
    LocalMux I__1695 (
            .O(N__8858),
            .I(N__8690));
    InMux I__1694 (
            .O(N__8857),
            .I(N__8681));
    InMux I__1693 (
            .O(N__8856),
            .I(N__8681));
    InMux I__1692 (
            .O(N__8855),
            .I(N__8681));
    InMux I__1691 (
            .O(N__8854),
            .I(N__8681));
    Span4Mux_v I__1690 (
            .O(N__8851),
            .I(N__8670));
    Span4Mux_h I__1689 (
            .O(N__8848),
            .I(N__8670));
    Span4Mux_v I__1688 (
            .O(N__8845),
            .I(N__8670));
    LocalMux I__1687 (
            .O(N__8834),
            .I(N__8670));
    LocalMux I__1686 (
            .O(N__8827),
            .I(N__8670));
    LocalMux I__1685 (
            .O(N__8824),
            .I(N__8657));
    LocalMux I__1684 (
            .O(N__8817),
            .I(N__8657));
    LocalMux I__1683 (
            .O(N__8804),
            .I(N__8657));
    LocalMux I__1682 (
            .O(N__8789),
            .I(N__8657));
    LocalMux I__1681 (
            .O(N__8778),
            .I(N__8657));
    LocalMux I__1680 (
            .O(N__8769),
            .I(N__8657));
    InMux I__1679 (
            .O(N__8768),
            .I(N__8654));
    LocalMux I__1678 (
            .O(N__8765),
            .I(N__8645));
    LocalMux I__1677 (
            .O(N__8756),
            .I(N__8645));
    Span4Mux_v I__1676 (
            .O(N__8751),
            .I(N__8640));
    LocalMux I__1675 (
            .O(N__8742),
            .I(N__8640));
    LocalMux I__1674 (
            .O(N__8725),
            .I(N__8637));
    InMux I__1673 (
            .O(N__8724),
            .I(N__8626));
    InMux I__1672 (
            .O(N__8723),
            .I(N__8626));
    InMux I__1671 (
            .O(N__8722),
            .I(N__8626));
    InMux I__1670 (
            .O(N__8721),
            .I(N__8626));
    InMux I__1669 (
            .O(N__8720),
            .I(N__8626));
    InMux I__1668 (
            .O(N__8719),
            .I(N__8611));
    InMux I__1667 (
            .O(N__8718),
            .I(N__8611));
    InMux I__1666 (
            .O(N__8717),
            .I(N__8611));
    InMux I__1665 (
            .O(N__8716),
            .I(N__8611));
    InMux I__1664 (
            .O(N__8715),
            .I(N__8611));
    InMux I__1663 (
            .O(N__8714),
            .I(N__8611));
    InMux I__1662 (
            .O(N__8713),
            .I(N__8611));
    InMux I__1661 (
            .O(N__8712),
            .I(N__8604));
    InMux I__1660 (
            .O(N__8711),
            .I(N__8604));
    InMux I__1659 (
            .O(N__8710),
            .I(N__8604));
    InMux I__1658 (
            .O(N__8709),
            .I(N__8601));
    Span4Mux_v I__1657 (
            .O(N__8698),
            .I(N__8592));
    Span4Mux_v I__1656 (
            .O(N__8695),
            .I(N__8592));
    Span4Mux_v I__1655 (
            .O(N__8690),
            .I(N__8592));
    LocalMux I__1654 (
            .O(N__8681),
            .I(N__8592));
    Span4Mux_h I__1653 (
            .O(N__8670),
            .I(N__8585));
    Span4Mux_v I__1652 (
            .O(N__8657),
            .I(N__8585));
    LocalMux I__1651 (
            .O(N__8654),
            .I(N__8585));
    InMux I__1650 (
            .O(N__8653),
            .I(N__8576));
    InMux I__1649 (
            .O(N__8652),
            .I(N__8576));
    InMux I__1648 (
            .O(N__8651),
            .I(N__8576));
    InMux I__1647 (
            .O(N__8650),
            .I(N__8576));
    Odrv12 I__1646 (
            .O(N__8645),
            .I(\FSM_TEST_inst_slow.current_stateZ1Z_0 ));
    Odrv4 I__1645 (
            .O(N__8640),
            .I(\FSM_TEST_inst_slow.current_stateZ1Z_0 ));
    Odrv4 I__1644 (
            .O(N__8637),
            .I(\FSM_TEST_inst_slow.current_stateZ1Z_0 ));
    LocalMux I__1643 (
            .O(N__8626),
            .I(\FSM_TEST_inst_slow.current_stateZ1Z_0 ));
    LocalMux I__1642 (
            .O(N__8611),
            .I(\FSM_TEST_inst_slow.current_stateZ1Z_0 ));
    LocalMux I__1641 (
            .O(N__8604),
            .I(\FSM_TEST_inst_slow.current_stateZ1Z_0 ));
    LocalMux I__1640 (
            .O(N__8601),
            .I(\FSM_TEST_inst_slow.current_stateZ1Z_0 ));
    Odrv4 I__1639 (
            .O(N__8592),
            .I(\FSM_TEST_inst_slow.current_stateZ1Z_0 ));
    Odrv4 I__1638 (
            .O(N__8585),
            .I(\FSM_TEST_inst_slow.current_stateZ1Z_0 ));
    LocalMux I__1637 (
            .O(N__8576),
            .I(\FSM_TEST_inst_slow.current_stateZ1Z_0 ));
    CascadeMux I__1636 (
            .O(N__8555),
            .I(N__8552));
    InMux I__1635 (
            .O(N__8552),
            .I(N__8549));
    LocalMux I__1634 (
            .O(N__8549),
            .I(counter_RNIFD27_2));
    InMux I__1633 (
            .O(N__8546),
            .I(N__8543));
    LocalMux I__1632 (
            .O(N__8543),
            .I(N__8540));
    Span4Mux_h I__1631 (
            .O(N__8540),
            .I(N__8537));
    Span4Mux_h I__1630 (
            .O(N__8537),
            .I(N__8530));
    InMux I__1629 (
            .O(N__8536),
            .I(N__8527));
    InMux I__1628 (
            .O(N__8535),
            .I(N__8520));
    InMux I__1627 (
            .O(N__8534),
            .I(N__8520));
    InMux I__1626 (
            .O(N__8533),
            .I(N__8520));
    Odrv4 I__1625 (
            .O(N__8530),
            .I(clk_continuous_slow));
    LocalMux I__1624 (
            .O(N__8527),
            .I(clk_continuous_slow));
    LocalMux I__1623 (
            .O(N__8520),
            .I(clk_continuous_slow));
    InMux I__1622 (
            .O(N__8513),
            .I(N__8509));
    InMux I__1621 (
            .O(N__8512),
            .I(N__8506));
    LocalMux I__1620 (
            .O(N__8509),
            .I(N__8503));
    LocalMux I__1619 (
            .O(N__8506),
            .I(\FSM_TEST_inst_slow.aux_selection_slow_0 ));
    Odrv4 I__1618 (
            .O(N__8503),
            .I(\FSM_TEST_inst_slow.aux_selection_slow_0 ));
    CascadeMux I__1617 (
            .O(N__8498),
            .I(N__8493));
    InMux I__1616 (
            .O(N__8497),
            .I(N__8490));
    InMux I__1615 (
            .O(N__8496),
            .I(N__8487));
    InMux I__1614 (
            .O(N__8493),
            .I(N__8483));
    LocalMux I__1613 (
            .O(N__8490),
            .I(N__8478));
    LocalMux I__1612 (
            .O(N__8487),
            .I(N__8478));
    InMux I__1611 (
            .O(N__8486),
            .I(N__8475));
    LocalMux I__1610 (
            .O(N__8483),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_fastZ0Z_1 ));
    Odrv4 I__1609 (
            .O(N__8478),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_fastZ0Z_1 ));
    LocalMux I__1608 (
            .O(N__8475),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_fastZ0Z_1 ));
    CascadeMux I__1607 (
            .O(N__8468),
            .I(N__8464));
    InMux I__1606 (
            .O(N__8467),
            .I(N__8457));
    InMux I__1605 (
            .O(N__8464),
            .I(N__8457));
    CascadeMux I__1604 (
            .O(N__8463),
            .I(N__8451));
    InMux I__1603 (
            .O(N__8462),
            .I(N__8447));
    LocalMux I__1602 (
            .O(N__8457),
            .I(N__8444));
    InMux I__1601 (
            .O(N__8456),
            .I(N__8441));
    InMux I__1600 (
            .O(N__8455),
            .I(N__8434));
    InMux I__1599 (
            .O(N__8454),
            .I(N__8434));
    InMux I__1598 (
            .O(N__8451),
            .I(N__8434));
    InMux I__1597 (
            .O(N__8450),
            .I(N__8429));
    LocalMux I__1596 (
            .O(N__8447),
            .I(N__8420));
    Span4Mux_v I__1595 (
            .O(N__8444),
            .I(N__8420));
    LocalMux I__1594 (
            .O(N__8441),
            .I(N__8420));
    LocalMux I__1593 (
            .O(N__8434),
            .I(N__8420));
    InMux I__1592 (
            .O(N__8433),
            .I(N__8415));
    InMux I__1591 (
            .O(N__8432),
            .I(N__8415));
    LocalMux I__1590 (
            .O(N__8429),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_1_repZ0Z1 ));
    Odrv4 I__1589 (
            .O(N__8420),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_1_repZ0Z1 ));
    LocalMux I__1588 (
            .O(N__8415),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_1_repZ0Z1 ));
    InMux I__1587 (
            .O(N__8408),
            .I(N__8405));
    LocalMux I__1586 (
            .O(N__8405),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_76 ));
    InMux I__1585 (
            .O(N__8402),
            .I(N__8399));
    LocalMux I__1584 (
            .O(N__8399),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_54 ));
    InMux I__1583 (
            .O(N__8396),
            .I(N__8393));
    LocalMux I__1582 (
            .O(N__8393),
            .I(\FSM_TEST_inst_RAPIDA.CLK_uC_2Z0Z_0 ));
    InMux I__1581 (
            .O(N__8390),
            .I(N__8387));
    LocalMux I__1580 (
            .O(N__8387),
            .I(\FSM_TEST_inst_RAPIDA.CLK_uC_6bZ0Z_0 ));
    CascadeMux I__1579 (
            .O(N__8384),
            .I(N__8380));
    InMux I__1578 (
            .O(N__8383),
            .I(N__8375));
    InMux I__1577 (
            .O(N__8380),
            .I(N__8375));
    LocalMux I__1576 (
            .O(N__8375),
            .I(\FSM_TEST_inst_RAPIDA.CLK_uCZ0 ));
    InMux I__1575 (
            .O(N__8372),
            .I(N__8369));
    LocalMux I__1574 (
            .O(N__8369),
            .I(\FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5DZ0Z1 ));
    InMux I__1573 (
            .O(N__8366),
            .I(N__8362));
    InMux I__1572 (
            .O(N__8365),
            .I(N__8359));
    LocalMux I__1571 (
            .O(N__8362),
            .I(N_3_0));
    LocalMux I__1570 (
            .O(N__8359),
            .I(N_3_0));
    InMux I__1569 (
            .O(N__8354),
            .I(N__8345));
    InMux I__1568 (
            .O(N__8353),
            .I(N__8345));
    InMux I__1567 (
            .O(N__8352),
            .I(N__8342));
    InMux I__1566 (
            .O(N__8351),
            .I(N__8339));
    InMux I__1565 (
            .O(N__8350),
            .I(N__8336));
    LocalMux I__1564 (
            .O(N__8345),
            .I(N_4_0));
    LocalMux I__1563 (
            .O(N__8342),
            .I(N_4_0));
    LocalMux I__1562 (
            .O(N__8339),
            .I(N_4_0));
    LocalMux I__1561 (
            .O(N__8336),
            .I(N_4_0));
    InMux I__1560 (
            .O(N__8327),
            .I(N__8323));
    CascadeMux I__1559 (
            .O(N__8326),
            .I(N__8320));
    LocalMux I__1558 (
            .O(N__8323),
            .I(N__8317));
    InMux I__1557 (
            .O(N__8320),
            .I(N__8314));
    Span4Mux_v I__1556 (
            .O(N__8317),
            .I(N__8309));
    LocalMux I__1555 (
            .O(N__8314),
            .I(N__8309));
    Span4Mux_h I__1554 (
            .O(N__8309),
            .I(N__8306));
    Odrv4 I__1553 (
            .O(N__8306),
            .I(CLK_uC_6c_0));
    IoInMux I__1552 (
            .O(N__8303),
            .I(N__8300));
    LocalMux I__1551 (
            .O(N__8300),
            .I(N__8297));
    Span4Mux_s1_v I__1550 (
            .O(N__8297),
            .I(N__8294));
    Span4Mux_v I__1549 (
            .O(N__8294),
            .I(N__8291));
    Sp12to4 I__1548 (
            .O(N__8291),
            .I(N__8287));
    InMux I__1547 (
            .O(N__8290),
            .I(N__8284));
    Span12Mux_h I__1546 (
            .O(N__8287),
            .I(N__8281));
    LocalMux I__1545 (
            .O(N__8284),
            .I(N__8278));
    Odrv12 I__1544 (
            .O(N__8281),
            .I(clk_output_c));
    Odrv4 I__1543 (
            .O(N__8278),
            .I(clk_output_c));
    InMux I__1542 (
            .O(N__8273),
            .I(N__8270));
    LocalMux I__1541 (
            .O(N__8270),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_6 ));
    InMux I__1540 (
            .O(N__8267),
            .I(N__8264));
    LocalMux I__1539 (
            .O(N__8264),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_7 ));
    InMux I__1538 (
            .O(N__8261),
            .I(N__8258));
    LocalMux I__1537 (
            .O(N__8258),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_8 ));
    InMux I__1536 (
            .O(N__8255),
            .I(N__8252));
    LocalMux I__1535 (
            .O(N__8252),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_9 ));
    InMux I__1534 (
            .O(N__8249),
            .I(N__8246));
    LocalMux I__1533 (
            .O(N__8246),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_11 ));
    InMux I__1532 (
            .O(N__8243),
            .I(N__8240));
    LocalMux I__1531 (
            .O(N__8240),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_12 ));
    CEMux I__1530 (
            .O(N__8237),
            .I(N__8234));
    LocalMux I__1529 (
            .O(N__8234),
            .I(N__8229));
    CEMux I__1528 (
            .O(N__8233),
            .I(N__8226));
    CEMux I__1527 (
            .O(N__8232),
            .I(N__8223));
    Span4Mux_h I__1526 (
            .O(N__8229),
            .I(N__8218));
    LocalMux I__1525 (
            .O(N__8226),
            .I(N__8218));
    LocalMux I__1524 (
            .O(N__8223),
            .I(N__8215));
    Odrv4 I__1523 (
            .O(N__8218),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_RNI78E11Z0Z_1 ));
    Odrv12 I__1522 (
            .O(N__8215),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_RNI78E11Z0Z_1 ));
    InMux I__1521 (
            .O(N__8210),
            .I(N__8207));
    LocalMux I__1520 (
            .O(N__8207),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_27 ));
    InMux I__1519 (
            .O(N__8204),
            .I(N__8201));
    LocalMux I__1518 (
            .O(N__8201),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_28 ));
    InMux I__1517 (
            .O(N__8198),
            .I(N__8195));
    LocalMux I__1516 (
            .O(N__8195),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_59 ));
    InMux I__1515 (
            .O(N__8192),
            .I(N__8186));
    InMux I__1514 (
            .O(N__8191),
            .I(N__8186));
    LocalMux I__1513 (
            .O(N__8186),
            .I(N__8183));
    Odrv4 I__1512 (
            .O(N__8183),
            .I(\FSM_TEST_inst_RAPIDA.N_101_0 ));
    CascadeMux I__1511 (
            .O(N__8180),
            .I(N__8176));
    InMux I__1510 (
            .O(N__8179),
            .I(N__8172));
    InMux I__1509 (
            .O(N__8176),
            .I(N__8169));
    InMux I__1508 (
            .O(N__8175),
            .I(N__8166));
    LocalMux I__1507 (
            .O(N__8172),
            .I(N__8163));
    LocalMux I__1506 (
            .O(N__8169),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_10 ));
    LocalMux I__1505 (
            .O(N__8166),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_10 ));
    Odrv4 I__1504 (
            .O(N__8163),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_10 ));
    InMux I__1503 (
            .O(N__8156),
            .I(N__8150));
    InMux I__1502 (
            .O(N__8155),
            .I(N__8150));
    LocalMux I__1501 (
            .O(N__8150),
            .I(N__8147));
    Span4Mux_v I__1500 (
            .O(N__8147),
            .I(N__8144));
    Span4Mux_h I__1499 (
            .O(N__8144),
            .I(N__8141));
    Sp12to4 I__1498 (
            .O(N__8141),
            .I(N__8138));
    Span12Mux_h I__1497 (
            .O(N__8138),
            .I(N__8135));
    Odrv12 I__1496 (
            .O(N__8135),
            .I(miso_input_c));
    InMux I__1495 (
            .O(N__8132),
            .I(N__8128));
    InMux I__1494 (
            .O(N__8131),
            .I(N__8125));
    LocalMux I__1493 (
            .O(N__8128),
            .I(N__8118));
    LocalMux I__1492 (
            .O(N__8125),
            .I(N__8118));
    InMux I__1491 (
            .O(N__8124),
            .I(N__8113));
    InMux I__1490 (
            .O(N__8123),
            .I(N__8113));
    Span4Mux_h I__1489 (
            .O(N__8118),
            .I(N__8110));
    LocalMux I__1488 (
            .O(N__8113),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_0 ));
    Odrv4 I__1487 (
            .O(N__8110),
            .I(\config_register_latched_dec_inst.DYNSRZ0Z_0 ));
    InMux I__1486 (
            .O(N__8105),
            .I(N__8102));
    LocalMux I__1485 (
            .O(N__8102),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_10 ));
    InMux I__1484 (
            .O(N__8099),
            .I(N__8096));
    LocalMux I__1483 (
            .O(N__8096),
            .I(N__8093));
    Span4Mux_h I__1482 (
            .O(N__8093),
            .I(N__8090));
    Odrv4 I__1481 (
            .O(N__8090),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_15 ));
    CascadeMux I__1480 (
            .O(N__8087),
            .I(clk_out_RNI3LEM_cascade_));
    CascadeMux I__1479 (
            .O(N__8084),
            .I(\FSM_TEST_inst_RAPIDA.N_100_li_cascade_ ));
    CascadeMux I__1478 (
            .O(N__8081),
            .I(\FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5DZ0Z1_cascade_ ));
    CEMux I__1477 (
            .O(N__8078),
            .I(N__8075));
    LocalMux I__1476 (
            .O(N__8075),
            .I(N__8072));
    Odrv4 I__1475 (
            .O(N__8072),
            .I(N_378_i));
    InMux I__1474 (
            .O(N__8069),
            .I(N__8063));
    InMux I__1473 (
            .O(N__8068),
            .I(N__8063));
    LocalMux I__1472 (
            .O(N__8063),
            .I(N__8058));
    InMux I__1471 (
            .O(N__8062),
            .I(N__8053));
    InMux I__1470 (
            .O(N__8061),
            .I(N__8053));
    Span4Mux_h I__1469 (
            .O(N__8058),
            .I(N__8050));
    LocalMux I__1468 (
            .O(N__8053),
            .I(flag_signal));
    Odrv4 I__1467 (
            .O(N__8050),
            .I(flag_signal));
    InMux I__1466 (
            .O(N__8045),
            .I(N__8042));
    LocalMux I__1465 (
            .O(N__8042),
            .I(mosi_fast));
    InMux I__1464 (
            .O(N__8039),
            .I(N__8036));
    LocalMux I__1463 (
            .O(N__8036),
            .I(N__8033));
    Span4Mux_h I__1462 (
            .O(N__8033),
            .I(N__8030));
    Odrv4 I__1461 (
            .O(N__8030),
            .I(mosi_slow));
    IoInMux I__1460 (
            .O(N__8027),
            .I(N__8024));
    LocalMux I__1459 (
            .O(N__8024),
            .I(N__8021));
    IoSpan4Mux I__1458 (
            .O(N__8021),
            .I(N__8018));
    Sp12to4 I__1457 (
            .O(N__8018),
            .I(N__8015));
    Span12Mux_s7_h I__1456 (
            .O(N__8015),
            .I(N__8012));
    Span12Mux_h I__1455 (
            .O(N__8012),
            .I(N__8009));
    Span12Mux_v I__1454 (
            .O(N__8009),
            .I(N__8006));
    Odrv12 I__1453 (
            .O(N__8006),
            .I(mosi_output_c));
    InMux I__1452 (
            .O(N__8003),
            .I(N__7999));
    CascadeMux I__1451 (
            .O(N__8002),
            .I(N__7996));
    LocalMux I__1450 (
            .O(N__7999),
            .I(N__7993));
    InMux I__1449 (
            .O(N__7996),
            .I(N__7990));
    Odrv4 I__1448 (
            .O(N__7993),
            .I(\config_register_latched_dec_inst.DYNCNF_1Z0Z_10 ));
    LocalMux I__1447 (
            .O(N__7990),
            .I(\config_register_latched_dec_inst.DYNCNF_1Z0Z_10 ));
    IoInMux I__1446 (
            .O(N__7985),
            .I(N__7982));
    LocalMux I__1445 (
            .O(N__7982),
            .I(N__7979));
    IoSpan4Mux I__1444 (
            .O(N__7979),
            .I(N__7976));
    Sp12to4 I__1443 (
            .O(N__7976),
            .I(N__7973));
    Span12Mux_h I__1442 (
            .O(N__7973),
            .I(N__7970));
    Odrv12 I__1441 (
            .O(N__7970),
            .I(s14_c));
    CEMux I__1440 (
            .O(N__7967),
            .I(N__7964));
    LocalMux I__1439 (
            .O(N__7964),
            .I(N__7961));
    Odrv12 I__1438 (
            .O(N__7961),
            .I(\config_register_latched_dec_inst.N_378_i_i ));
    InMux I__1437 (
            .O(N__7958),
            .I(N__7955));
    LocalMux I__1436 (
            .O(N__7955),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_64 ));
    InMux I__1435 (
            .O(N__7952),
            .I(N__7949));
    LocalMux I__1434 (
            .O(N__7949),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_65 ));
    InMux I__1433 (
            .O(N__7946),
            .I(N__7943));
    LocalMux I__1432 (
            .O(N__7943),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_62 ));
    CascadeMux I__1431 (
            .O(N__7940),
            .I(N__7935));
    CascadeMux I__1430 (
            .O(N__7939),
            .I(N__7932));
    CascadeMux I__1429 (
            .O(N__7938),
            .I(N__7910));
    InMux I__1428 (
            .O(N__7935),
            .I(N__7892));
    InMux I__1427 (
            .O(N__7932),
            .I(N__7892));
    InMux I__1426 (
            .O(N__7931),
            .I(N__7892));
    InMux I__1425 (
            .O(N__7930),
            .I(N__7889));
    InMux I__1424 (
            .O(N__7929),
            .I(N__7882));
    CascadeMux I__1423 (
            .O(N__7928),
            .I(N__7872));
    CascadeMux I__1422 (
            .O(N__7927),
            .I(N__7869));
    CascadeMux I__1421 (
            .O(N__7926),
            .I(N__7866));
    CascadeMux I__1420 (
            .O(N__7925),
            .I(N__7860));
    CascadeMux I__1419 (
            .O(N__7924),
            .I(N__7855));
    CascadeMux I__1418 (
            .O(N__7923),
            .I(N__7852));
    CascadeMux I__1417 (
            .O(N__7922),
            .I(N__7845));
    CascadeMux I__1416 (
            .O(N__7921),
            .I(N__7842));
    CascadeMux I__1415 (
            .O(N__7920),
            .I(N__7838));
    InMux I__1414 (
            .O(N__7919),
            .I(N__7824));
    CascadeMux I__1413 (
            .O(N__7918),
            .I(N__7821));
    CascadeMux I__1412 (
            .O(N__7917),
            .I(N__7818));
    CascadeMux I__1411 (
            .O(N__7916),
            .I(N__7815));
    CascadeMux I__1410 (
            .O(N__7915),
            .I(N__7808));
    CascadeMux I__1409 (
            .O(N__7914),
            .I(N__7804));
    CascadeMux I__1408 (
            .O(N__7913),
            .I(N__7801));
    InMux I__1407 (
            .O(N__7910),
            .I(N__7791));
    InMux I__1406 (
            .O(N__7909),
            .I(N__7791));
    InMux I__1405 (
            .O(N__7908),
            .I(N__7786));
    InMux I__1404 (
            .O(N__7907),
            .I(N__7786));
    CascadeMux I__1403 (
            .O(N__7906),
            .I(N__7782));
    CascadeMux I__1402 (
            .O(N__7905),
            .I(N__7778));
    CascadeMux I__1401 (
            .O(N__7904),
            .I(N__7775));
    CascadeMux I__1400 (
            .O(N__7903),
            .I(N__7770));
    CascadeMux I__1399 (
            .O(N__7902),
            .I(N__7767));
    CascadeMux I__1398 (
            .O(N__7901),
            .I(N__7763));
    CascadeMux I__1397 (
            .O(N__7900),
            .I(N__7758));
    CascadeMux I__1396 (
            .O(N__7899),
            .I(N__7754));
    LocalMux I__1395 (
            .O(N__7892),
            .I(N__7749));
    LocalMux I__1394 (
            .O(N__7889),
            .I(N__7746));
    InMux I__1393 (
            .O(N__7888),
            .I(N__7743));
    InMux I__1392 (
            .O(N__7887),
            .I(N__7736));
    InMux I__1391 (
            .O(N__7886),
            .I(N__7736));
    InMux I__1390 (
            .O(N__7885),
            .I(N__7736));
    LocalMux I__1389 (
            .O(N__7882),
            .I(N__7733));
    InMux I__1388 (
            .O(N__7881),
            .I(N__7722));
    InMux I__1387 (
            .O(N__7880),
            .I(N__7722));
    InMux I__1386 (
            .O(N__7879),
            .I(N__7722));
    InMux I__1385 (
            .O(N__7878),
            .I(N__7722));
    InMux I__1384 (
            .O(N__7877),
            .I(N__7722));
    InMux I__1383 (
            .O(N__7876),
            .I(N__7707));
    InMux I__1382 (
            .O(N__7875),
            .I(N__7707));
    InMux I__1381 (
            .O(N__7872),
            .I(N__7707));
    InMux I__1380 (
            .O(N__7869),
            .I(N__7707));
    InMux I__1379 (
            .O(N__7866),
            .I(N__7707));
    InMux I__1378 (
            .O(N__7865),
            .I(N__7707));
    InMux I__1377 (
            .O(N__7864),
            .I(N__7707));
    InMux I__1376 (
            .O(N__7863),
            .I(N__7700));
    InMux I__1375 (
            .O(N__7860),
            .I(N__7700));
    InMux I__1374 (
            .O(N__7859),
            .I(N__7700));
    InMux I__1373 (
            .O(N__7858),
            .I(N__7691));
    InMux I__1372 (
            .O(N__7855),
            .I(N__7691));
    InMux I__1371 (
            .O(N__7852),
            .I(N__7691));
    InMux I__1370 (
            .O(N__7851),
            .I(N__7691));
    InMux I__1369 (
            .O(N__7850),
            .I(N__7688));
    InMux I__1368 (
            .O(N__7849),
            .I(N__7685));
    InMux I__1367 (
            .O(N__7848),
            .I(N__7682));
    InMux I__1366 (
            .O(N__7845),
            .I(N__7671));
    InMux I__1365 (
            .O(N__7842),
            .I(N__7671));
    InMux I__1364 (
            .O(N__7841),
            .I(N__7671));
    InMux I__1363 (
            .O(N__7838),
            .I(N__7671));
    InMux I__1362 (
            .O(N__7837),
            .I(N__7671));
    InMux I__1361 (
            .O(N__7836),
            .I(N__7654));
    InMux I__1360 (
            .O(N__7835),
            .I(N__7654));
    InMux I__1359 (
            .O(N__7834),
            .I(N__7654));
    InMux I__1358 (
            .O(N__7833),
            .I(N__7654));
    InMux I__1357 (
            .O(N__7832),
            .I(N__7645));
    InMux I__1356 (
            .O(N__7831),
            .I(N__7645));
    InMux I__1355 (
            .O(N__7830),
            .I(N__7645));
    InMux I__1354 (
            .O(N__7829),
            .I(N__7645));
    CascadeMux I__1353 (
            .O(N__7828),
            .I(N__7641));
    InMux I__1352 (
            .O(N__7827),
            .I(N__7635));
    LocalMux I__1351 (
            .O(N__7824),
            .I(N__7632));
    InMux I__1350 (
            .O(N__7821),
            .I(N__7621));
    InMux I__1349 (
            .O(N__7818),
            .I(N__7621));
    InMux I__1348 (
            .O(N__7815),
            .I(N__7621));
    InMux I__1347 (
            .O(N__7814),
            .I(N__7621));
    InMux I__1346 (
            .O(N__7813),
            .I(N__7621));
    InMux I__1345 (
            .O(N__7812),
            .I(N__7617));
    InMux I__1344 (
            .O(N__7811),
            .I(N__7614));
    InMux I__1343 (
            .O(N__7808),
            .I(N__7609));
    InMux I__1342 (
            .O(N__7807),
            .I(N__7609));
    InMux I__1341 (
            .O(N__7804),
            .I(N__7602));
    InMux I__1340 (
            .O(N__7801),
            .I(N__7602));
    InMux I__1339 (
            .O(N__7800),
            .I(N__7602));
    InMux I__1338 (
            .O(N__7799),
            .I(N__7593));
    InMux I__1337 (
            .O(N__7798),
            .I(N__7593));
    InMux I__1336 (
            .O(N__7797),
            .I(N__7593));
    InMux I__1335 (
            .O(N__7796),
            .I(N__7593));
    LocalMux I__1334 (
            .O(N__7791),
            .I(N__7588));
    LocalMux I__1333 (
            .O(N__7786),
            .I(N__7588));
    InMux I__1332 (
            .O(N__7785),
            .I(N__7573));
    InMux I__1331 (
            .O(N__7782),
            .I(N__7573));
    InMux I__1330 (
            .O(N__7781),
            .I(N__7573));
    InMux I__1329 (
            .O(N__7778),
            .I(N__7573));
    InMux I__1328 (
            .O(N__7775),
            .I(N__7573));
    InMux I__1327 (
            .O(N__7774),
            .I(N__7573));
    InMux I__1326 (
            .O(N__7773),
            .I(N__7573));
    InMux I__1325 (
            .O(N__7770),
            .I(N__7548));
    InMux I__1324 (
            .O(N__7767),
            .I(N__7548));
    InMux I__1323 (
            .O(N__7766),
            .I(N__7548));
    InMux I__1322 (
            .O(N__7763),
            .I(N__7548));
    InMux I__1321 (
            .O(N__7762),
            .I(N__7548));
    InMux I__1320 (
            .O(N__7761),
            .I(N__7548));
    InMux I__1319 (
            .O(N__7758),
            .I(N__7537));
    InMux I__1318 (
            .O(N__7757),
            .I(N__7537));
    InMux I__1317 (
            .O(N__7754),
            .I(N__7537));
    InMux I__1316 (
            .O(N__7753),
            .I(N__7537));
    InMux I__1315 (
            .O(N__7752),
            .I(N__7537));
    Span4Mux_v I__1314 (
            .O(N__7749),
            .I(N__7525));
    Span4Mux_v I__1313 (
            .O(N__7746),
            .I(N__7525));
    LocalMux I__1312 (
            .O(N__7743),
            .I(N__7525));
    LocalMux I__1311 (
            .O(N__7736),
            .I(N__7525));
    Span4Mux_v I__1310 (
            .O(N__7733),
            .I(N__7514));
    LocalMux I__1309 (
            .O(N__7722),
            .I(N__7514));
    LocalMux I__1308 (
            .O(N__7707),
            .I(N__7514));
    LocalMux I__1307 (
            .O(N__7700),
            .I(N__7514));
    LocalMux I__1306 (
            .O(N__7691),
            .I(N__7514));
    LocalMux I__1305 (
            .O(N__7688),
            .I(N__7509));
    LocalMux I__1304 (
            .O(N__7685),
            .I(N__7509));
    LocalMux I__1303 (
            .O(N__7682),
            .I(N__7504));
    LocalMux I__1302 (
            .O(N__7671),
            .I(N__7504));
    InMux I__1301 (
            .O(N__7670),
            .I(N__7487));
    InMux I__1300 (
            .O(N__7669),
            .I(N__7487));
    InMux I__1299 (
            .O(N__7668),
            .I(N__7487));
    InMux I__1298 (
            .O(N__7667),
            .I(N__7487));
    InMux I__1297 (
            .O(N__7666),
            .I(N__7487));
    InMux I__1296 (
            .O(N__7665),
            .I(N__7487));
    InMux I__1295 (
            .O(N__7664),
            .I(N__7487));
    InMux I__1294 (
            .O(N__7663),
            .I(N__7487));
    LocalMux I__1293 (
            .O(N__7654),
            .I(N__7482));
    LocalMux I__1292 (
            .O(N__7645),
            .I(N__7482));
    InMux I__1291 (
            .O(N__7644),
            .I(N__7471));
    InMux I__1290 (
            .O(N__7641),
            .I(N__7471));
    InMux I__1289 (
            .O(N__7640),
            .I(N__7471));
    InMux I__1288 (
            .O(N__7639),
            .I(N__7471));
    InMux I__1287 (
            .O(N__7638),
            .I(N__7471));
    LocalMux I__1286 (
            .O(N__7635),
            .I(N__7468));
    Span4Mux_h I__1285 (
            .O(N__7632),
            .I(N__7463));
    LocalMux I__1284 (
            .O(N__7621),
            .I(N__7463));
    InMux I__1283 (
            .O(N__7620),
            .I(N__7460));
    LocalMux I__1282 (
            .O(N__7617),
            .I(N__7454));
    LocalMux I__1281 (
            .O(N__7614),
            .I(N__7447));
    LocalMux I__1280 (
            .O(N__7609),
            .I(N__7447));
    LocalMux I__1279 (
            .O(N__7602),
            .I(N__7447));
    LocalMux I__1278 (
            .O(N__7593),
            .I(N__7444));
    Span4Mux_h I__1277 (
            .O(N__7588),
            .I(N__7439));
    LocalMux I__1276 (
            .O(N__7573),
            .I(N__7439));
    InMux I__1275 (
            .O(N__7572),
            .I(N__7432));
    InMux I__1274 (
            .O(N__7571),
            .I(N__7432));
    InMux I__1273 (
            .O(N__7570),
            .I(N__7432));
    InMux I__1272 (
            .O(N__7569),
            .I(N__7427));
    InMux I__1271 (
            .O(N__7568),
            .I(N__7427));
    InMux I__1270 (
            .O(N__7567),
            .I(N__7420));
    InMux I__1269 (
            .O(N__7566),
            .I(N__7420));
    InMux I__1268 (
            .O(N__7565),
            .I(N__7420));
    InMux I__1267 (
            .O(N__7564),
            .I(N__7411));
    InMux I__1266 (
            .O(N__7563),
            .I(N__7411));
    InMux I__1265 (
            .O(N__7562),
            .I(N__7411));
    InMux I__1264 (
            .O(N__7561),
            .I(N__7411));
    LocalMux I__1263 (
            .O(N__7548),
            .I(N__7406));
    LocalMux I__1262 (
            .O(N__7537),
            .I(N__7406));
    InMux I__1261 (
            .O(N__7536),
            .I(N__7399));
    InMux I__1260 (
            .O(N__7535),
            .I(N__7399));
    InMux I__1259 (
            .O(N__7534),
            .I(N__7399));
    Span4Mux_h I__1258 (
            .O(N__7525),
            .I(N__7392));
    Span4Mux_v I__1257 (
            .O(N__7514),
            .I(N__7392));
    Span4Mux_v I__1256 (
            .O(N__7509),
            .I(N__7392));
    Span4Mux_v I__1255 (
            .O(N__7504),
            .I(N__7383));
    LocalMux I__1254 (
            .O(N__7487),
            .I(N__7383));
    Span4Mux_v I__1253 (
            .O(N__7482),
            .I(N__7383));
    LocalMux I__1252 (
            .O(N__7471),
            .I(N__7383));
    Span4Mux_v I__1251 (
            .O(N__7468),
            .I(N__7376));
    Span4Mux_h I__1250 (
            .O(N__7463),
            .I(N__7376));
    LocalMux I__1249 (
            .O(N__7460),
            .I(N__7376));
    InMux I__1248 (
            .O(N__7459),
            .I(N__7369));
    InMux I__1247 (
            .O(N__7458),
            .I(N__7369));
    InMux I__1246 (
            .O(N__7457),
            .I(N__7369));
    Odrv12 I__1245 (
            .O(N__7454),
            .I(\FSM_TEST_inst_slow.current_stateZ0Z_1 ));
    Odrv12 I__1244 (
            .O(N__7447),
            .I(\FSM_TEST_inst_slow.current_stateZ0Z_1 ));
    Odrv4 I__1243 (
            .O(N__7444),
            .I(\FSM_TEST_inst_slow.current_stateZ0Z_1 ));
    Odrv4 I__1242 (
            .O(N__7439),
            .I(\FSM_TEST_inst_slow.current_stateZ0Z_1 ));
    LocalMux I__1241 (
            .O(N__7432),
            .I(\FSM_TEST_inst_slow.current_stateZ0Z_1 ));
    LocalMux I__1240 (
            .O(N__7427),
            .I(\FSM_TEST_inst_slow.current_stateZ0Z_1 ));
    LocalMux I__1239 (
            .O(N__7420),
            .I(\FSM_TEST_inst_slow.current_stateZ0Z_1 ));
    LocalMux I__1238 (
            .O(N__7411),
            .I(\FSM_TEST_inst_slow.current_stateZ0Z_1 ));
    Odrv4 I__1237 (
            .O(N__7406),
            .I(\FSM_TEST_inst_slow.current_stateZ0Z_1 ));
    LocalMux I__1236 (
            .O(N__7399),
            .I(\FSM_TEST_inst_slow.current_stateZ0Z_1 ));
    Odrv4 I__1235 (
            .O(N__7392),
            .I(\FSM_TEST_inst_slow.current_stateZ0Z_1 ));
    Odrv4 I__1234 (
            .O(N__7383),
            .I(\FSM_TEST_inst_slow.current_stateZ0Z_1 ));
    Odrv4 I__1233 (
            .O(N__7376),
            .I(\FSM_TEST_inst_slow.current_stateZ0Z_1 ));
    LocalMux I__1232 (
            .O(N__7369),
            .I(\FSM_TEST_inst_slow.current_stateZ0Z_1 ));
    InMux I__1231 (
            .O(N__7340),
            .I(N__7337));
    LocalMux I__1230 (
            .O(N__7337),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_63 ));
    CEMux I__1229 (
            .O(N__7334),
            .I(N__7259));
    CEMux I__1228 (
            .O(N__7333),
            .I(N__7259));
    CEMux I__1227 (
            .O(N__7332),
            .I(N__7259));
    CEMux I__1226 (
            .O(N__7331),
            .I(N__7259));
    CEMux I__1225 (
            .O(N__7330),
            .I(N__7259));
    CEMux I__1224 (
            .O(N__7329),
            .I(N__7259));
    CEMux I__1223 (
            .O(N__7328),
            .I(N__7259));
    CEMux I__1222 (
            .O(N__7327),
            .I(N__7259));
    CEMux I__1221 (
            .O(N__7326),
            .I(N__7259));
    CEMux I__1220 (
            .O(N__7325),
            .I(N__7259));
    CEMux I__1219 (
            .O(N__7324),
            .I(N__7259));
    CEMux I__1218 (
            .O(N__7323),
            .I(N__7259));
    CEMux I__1217 (
            .O(N__7322),
            .I(N__7259));
    CEMux I__1216 (
            .O(N__7321),
            .I(N__7259));
    CEMux I__1215 (
            .O(N__7320),
            .I(N__7259));
    CEMux I__1214 (
            .O(N__7319),
            .I(N__7259));
    CEMux I__1213 (
            .O(N__7318),
            .I(N__7259));
    CEMux I__1212 (
            .O(N__7317),
            .I(N__7259));
    CEMux I__1211 (
            .O(N__7316),
            .I(N__7259));
    CEMux I__1210 (
            .O(N__7315),
            .I(N__7259));
    CEMux I__1209 (
            .O(N__7314),
            .I(N__7259));
    CEMux I__1208 (
            .O(N__7313),
            .I(N__7259));
    CEMux I__1207 (
            .O(N__7312),
            .I(N__7259));
    CEMux I__1206 (
            .O(N__7311),
            .I(N__7259));
    CEMux I__1205 (
            .O(N__7310),
            .I(N__7259));
    GlobalMux I__1204 (
            .O(N__7259),
            .I(N__7256));
    gio2CtrlBuf I__1203 (
            .O(N__7256),
            .I(\FSM_TEST_inst_slow.N_374_g ));
    CascadeMux I__1202 (
            .O(N__7253),
            .I(counter_RNIFD27_2_cascade_));
    CascadeMux I__1201 (
            .O(N__7250),
            .I(N_3_0_cascade_));
    InMux I__1200 (
            .O(N__7247),
            .I(N__7244));
    LocalMux I__1199 (
            .O(N__7244),
            .I(N_2_0));
    CEMux I__1198 (
            .O(N__7241),
            .I(N__7235));
    InMux I__1197 (
            .O(N__7240),
            .I(N__7228));
    InMux I__1196 (
            .O(N__7239),
            .I(N__7228));
    InMux I__1195 (
            .O(N__7238),
            .I(N__7228));
    LocalMux I__1194 (
            .O(N__7235),
            .I(N__7222));
    LocalMux I__1193 (
            .O(N__7228),
            .I(N__7219));
    InMux I__1192 (
            .O(N__7227),
            .I(N__7212));
    InMux I__1191 (
            .O(N__7226),
            .I(N__7212));
    InMux I__1190 (
            .O(N__7225),
            .I(N__7212));
    Span4Mux_h I__1189 (
            .O(N__7222),
            .I(N__7205));
    Span4Mux_v I__1188 (
            .O(N__7219),
            .I(N__7200));
    LocalMux I__1187 (
            .O(N__7212),
            .I(N__7200));
    InMux I__1186 (
            .O(N__7211),
            .I(N__7191));
    InMux I__1185 (
            .O(N__7210),
            .I(N__7191));
    InMux I__1184 (
            .O(N__7209),
            .I(N__7191));
    InMux I__1183 (
            .O(N__7208),
            .I(N__7191));
    Odrv4 I__1182 (
            .O(N__7205),
            .I(counter_RNISR1F_2));
    Odrv4 I__1181 (
            .O(N__7200),
            .I(counter_RNISR1F_2));
    LocalMux I__1180 (
            .O(N__7191),
            .I(counter_RNISR1F_2));
    InMux I__1179 (
            .O(N__7184),
            .I(N__7181));
    LocalMux I__1178 (
            .O(N__7181),
            .I(\FSM_TEST_inst_RAPIDA.CLK_uC_3Z0Z_0 ));
    InMux I__1177 (
            .O(N__7178),
            .I(N__7175));
    LocalMux I__1176 (
            .O(N__7175),
            .I(\FSM_TEST_inst_RAPIDA.CLK_uC_4Z0Z_0 ));
    InMux I__1175 (
            .O(N__7172),
            .I(N__7169));
    LocalMux I__1174 (
            .O(N__7169),
            .I(\FSM_TEST_inst_RAPIDA.CLK_uC_5Z0Z_0 ));
    InMux I__1173 (
            .O(N__7166),
            .I(N__7163));
    LocalMux I__1172 (
            .O(N__7163),
            .I(\FSM_TEST_inst_RAPIDA.CLK_uC_6Z0Z_0 ));
    InMux I__1171 (
            .O(N__7160),
            .I(N__7157));
    LocalMux I__1170 (
            .O(N__7157),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_57 ));
    InMux I__1169 (
            .O(N__7154),
            .I(N__7151));
    LocalMux I__1168 (
            .O(N__7151),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_60 ));
    InMux I__1167 (
            .O(N__7148),
            .I(N__7145));
    LocalMux I__1166 (
            .O(N__7145),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_58 ));
    InMux I__1165 (
            .O(N__7142),
            .I(N__7139));
    LocalMux I__1164 (
            .O(N__7139),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_59 ));
    InMux I__1163 (
            .O(N__7136),
            .I(N__7133));
    LocalMux I__1162 (
            .O(N__7133),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_61 ));
    InMux I__1161 (
            .O(N__7130),
            .I(N__7127));
    LocalMux I__1160 (
            .O(N__7127),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_66 ));
    InMux I__1159 (
            .O(N__7124),
            .I(N__7121));
    LocalMux I__1158 (
            .O(N__7121),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_13 ));
    InMux I__1157 (
            .O(N__7118),
            .I(N__7115));
    LocalMux I__1156 (
            .O(N__7115),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_14 ));
    InMux I__1155 (
            .O(N__7112),
            .I(N__7109));
    LocalMux I__1154 (
            .O(N__7109),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_18 ));
    InMux I__1153 (
            .O(N__7106),
            .I(N__7103));
    LocalMux I__1152 (
            .O(N__7103),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_24 ));
    InMux I__1151 (
            .O(N__7100),
            .I(N__7097));
    LocalMux I__1150 (
            .O(N__7097),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_78 ));
    InMux I__1149 (
            .O(N__7094),
            .I(N__7091));
    LocalMux I__1148 (
            .O(N__7091),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_77 ));
    InMux I__1147 (
            .O(N__7088),
            .I(N__7085));
    LocalMux I__1146 (
            .O(N__7085),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_25 ));
    InMux I__1145 (
            .O(N__7082),
            .I(N__7079));
    LocalMux I__1144 (
            .O(N__7079),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_26 ));
    InMux I__1143 (
            .O(N__7076),
            .I(N__7073));
    LocalMux I__1142 (
            .O(N__7073),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_0 ));
    InMux I__1141 (
            .O(N__7070),
            .I(N__7067));
    LocalMux I__1140 (
            .O(N__7067),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_1 ));
    InMux I__1139 (
            .O(N__7064),
            .I(N__7061));
    LocalMux I__1138 (
            .O(N__7061),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_4 ));
    InMux I__1137 (
            .O(N__7058),
            .I(N__7055));
    LocalMux I__1136 (
            .O(N__7055),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_5 ));
    InMux I__1135 (
            .O(N__7052),
            .I(N__7049));
    LocalMux I__1134 (
            .O(N__7049),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_2 ));
    InMux I__1133 (
            .O(N__7046),
            .I(N__7043));
    LocalMux I__1132 (
            .O(N__7043),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_3 ));
    CascadeMux I__1131 (
            .O(N__7040),
            .I(\FSM_TEST_inst_RAPIDA.counter_din_3_i_0_2_cascade_ ));
    CascadeMux I__1130 (
            .O(N__7037),
            .I(\FSM_TEST_inst_RAPIDA.G_24_0_o4_2_cascade_ ));
    InMux I__1129 (
            .O(N__7034),
            .I(N__7031));
    LocalMux I__1128 (
            .O(N__7031),
            .I(N__7028));
    Odrv4 I__1127 (
            .O(N__7028),
            .I(\FSM_TEST_inst_RAPIDA.G_24_0_a4_0_1 ));
    CascadeMux I__1126 (
            .O(N__7025),
            .I(N__7022));
    InMux I__1125 (
            .O(N__7022),
            .I(N__7018));
    CascadeMux I__1124 (
            .O(N__7021),
            .I(N__7014));
    LocalMux I__1123 (
            .O(N__7018),
            .I(N__7011));
    CascadeMux I__1122 (
            .O(N__7017),
            .I(N__7008));
    InMux I__1121 (
            .O(N__7014),
            .I(N__7005));
    Span4Mux_h I__1120 (
            .O(N__7011),
            .I(N__7002));
    InMux I__1119 (
            .O(N__7008),
            .I(N__6999));
    LocalMux I__1118 (
            .O(N__7005),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_6 ));
    Odrv4 I__1117 (
            .O(N__7002),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_6 ));
    LocalMux I__1116 (
            .O(N__6999),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_6 ));
    InMux I__1115 (
            .O(N__6992),
            .I(N__6989));
    LocalMux I__1114 (
            .O(N__6989),
            .I(N__6986));
    Span4Mux_h I__1113 (
            .O(N__6986),
            .I(N__6980));
    InMux I__1112 (
            .O(N__6985),
            .I(N__6977));
    InMux I__1111 (
            .O(N__6984),
            .I(N__6972));
    InMux I__1110 (
            .O(N__6983),
            .I(N__6972));
    Odrv4 I__1109 (
            .O(N__6980),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_3 ));
    LocalMux I__1108 (
            .O(N__6977),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_3 ));
    LocalMux I__1107 (
            .O(N__6972),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_3 ));
    InMux I__1106 (
            .O(N__6965),
            .I(N__6962));
    LocalMux I__1105 (
            .O(N__6962),
            .I(\FSM_TEST_inst_RAPIDA.G_24_0_a4_0_5 ));
    InMux I__1104 (
            .O(N__6959),
            .I(N__6956));
    LocalMux I__1103 (
            .O(N__6956),
            .I(\FSM_TEST_inst_RAPIDA.N_18_0 ));
    CascadeMux I__1102 (
            .O(N__6953),
            .I(\FSM_TEST_inst_RAPIDA.G_24_0_a4_0_6_cascade_ ));
    InMux I__1101 (
            .O(N__6950),
            .I(N__6947));
    LocalMux I__1100 (
            .O(N__6947),
            .I(\FSM_TEST_inst_RAPIDA.N_9_1 ));
    InMux I__1099 (
            .O(N__6944),
            .I(N__6937));
    InMux I__1098 (
            .O(N__6943),
            .I(N__6937));
    CascadeMux I__1097 (
            .O(N__6942),
            .I(N__6934));
    LocalMux I__1096 (
            .O(N__6937),
            .I(N__6931));
    InMux I__1095 (
            .O(N__6934),
            .I(N__6928));
    Span4Mux_v I__1094 (
            .O(N__6931),
            .I(N__6925));
    LocalMux I__1093 (
            .O(N__6928),
            .I(\FSM_TEST_inst_slow.counter_dinZ0Z_3 ));
    Odrv4 I__1092 (
            .O(N__6925),
            .I(\FSM_TEST_inst_slow.counter_dinZ0Z_3 ));
    InMux I__1091 (
            .O(N__6920),
            .I(N__6917));
    LocalMux I__1090 (
            .O(N__6917),
            .I(N__6913));
    CascadeMux I__1089 (
            .O(N__6916),
            .I(N__6909));
    Span4Mux_h I__1088 (
            .O(N__6913),
            .I(N__6905));
    InMux I__1087 (
            .O(N__6912),
            .I(N__6898));
    InMux I__1086 (
            .O(N__6909),
            .I(N__6898));
    InMux I__1085 (
            .O(N__6908),
            .I(N__6898));
    Odrv4 I__1084 (
            .O(N__6905),
            .I(\FSM_TEST_inst_slow.counter_dinZ0Z_2 ));
    LocalMux I__1083 (
            .O(N__6898),
            .I(\FSM_TEST_inst_slow.counter_dinZ0Z_2 ));
    InMux I__1082 (
            .O(N__6893),
            .I(N__6884));
    InMux I__1081 (
            .O(N__6892),
            .I(N__6884));
    InMux I__1080 (
            .O(N__6891),
            .I(N__6884));
    LocalMux I__1079 (
            .O(N__6884),
            .I(N__6881));
    Span4Mux_v I__1078 (
            .O(N__6881),
            .I(N__6878));
    Odrv4 I__1077 (
            .O(N__6878),
            .I(\FSM_TEST_inst_slow.N_106_0 ));
    CascadeMux I__1076 (
            .O(N__6875),
            .I(\FSM_TEST_inst_slow.current_state_RNO_8Z0Z_0_cascade_ ));
    InMux I__1075 (
            .O(N__6872),
            .I(N__6869));
    LocalMux I__1074 (
            .O(N__6869),
            .I(\FSM_TEST_inst_slow.current_state_RNO_1Z0Z_0 ));
    InMux I__1073 (
            .O(N__6866),
            .I(N__6863));
    LocalMux I__1072 (
            .O(N__6863),
            .I(N__6860));
    Odrv4 I__1071 (
            .O(N__6860),
            .I(\FSM_TEST_inst_slow.N_134 ));
    CascadeMux I__1070 (
            .O(N__6857),
            .I(\FSM_TEST_inst_slow.current_state_RNO_2Z0Z_0_cascade_ ));
    IoInMux I__1069 (
            .O(N__6854),
            .I(N__6851));
    LocalMux I__1068 (
            .O(N__6851),
            .I(N__6848));
    Span4Mux_s1_v I__1067 (
            .O(N__6848),
            .I(N__6845));
    Sp12to4 I__1066 (
            .O(N__6845),
            .I(N__6842));
    Span12Mux_s11_h I__1065 (
            .O(N__6842),
            .I(N__6839));
    Span12Mux_v I__1064 (
            .O(N__6839),
            .I(N__6836));
    Odrv12 I__1063 (
            .O(N__6836),
            .I(s12_c));
    CascadeMux I__1062 (
            .O(N__6833),
            .I(N__6829));
    InMux I__1061 (
            .O(N__6832),
            .I(N__6824));
    InMux I__1060 (
            .O(N__6829),
            .I(N__6824));
    LocalMux I__1059 (
            .O(N__6824),
            .I(\config_register_latched_dec_inst.DYNCNF_1Z0Z_8 ));
    InMux I__1058 (
            .O(N__6821),
            .I(N__6815));
    InMux I__1057 (
            .O(N__6820),
            .I(N__6815));
    LocalMux I__1056 (
            .O(N__6815),
            .I(\config_register_latched_dec_inst.DYNCNF_1Z0Z_9 ));
    IoInMux I__1055 (
            .O(N__6812),
            .I(N__6809));
    LocalMux I__1054 (
            .O(N__6809),
            .I(N__6806));
    Span12Mux_s11_h I__1053 (
            .O(N__6806),
            .I(N__6803));
    Odrv12 I__1052 (
            .O(N__6803),
            .I(s13_c));
    InMux I__1051 (
            .O(N__6800),
            .I(N__6794));
    InMux I__1050 (
            .O(N__6799),
            .I(N__6794));
    LocalMux I__1049 (
            .O(N__6794),
            .I(\config_register_latched_dec_inst.DYNCNF_1Z0Z_0 ));
    InMux I__1048 (
            .O(N__6791),
            .I(N__6788));
    LocalMux I__1047 (
            .O(N__6788),
            .I(N__6785));
    Span4Mux_h I__1046 (
            .O(N__6785),
            .I(N__6782));
    Span4Mux_v I__1045 (
            .O(N__6782),
            .I(N__6779));
    Sp12to4 I__1044 (
            .O(N__6779),
            .I(N__6776));
    Span12Mux_v I__1043 (
            .O(N__6776),
            .I(N__6773));
    Odrv12 I__1042 (
            .O(N__6773),
            .I(\config_register_latched_dec_inst.DYNCNF_0 ));
    InMux I__1041 (
            .O(N__6770),
            .I(N__6767));
    LocalMux I__1040 (
            .O(N__6767),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_6 ));
    InMux I__1039 (
            .O(N__6764),
            .I(N__6761));
    LocalMux I__1038 (
            .O(N__6761),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_56 ));
    InMux I__1037 (
            .O(N__6758),
            .I(N__6755));
    LocalMux I__1036 (
            .O(N__6755),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_69 ));
    InMux I__1035 (
            .O(N__6752),
            .I(N__6749));
    LocalMux I__1034 (
            .O(N__6749),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_68 ));
    InMux I__1033 (
            .O(N__6746),
            .I(N__6743));
    LocalMux I__1032 (
            .O(N__6743),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_67 ));
    CascadeMux I__1031 (
            .O(N__6740),
            .I(\FSM_TEST_inst_slow.N_108_li_cascade_ ));
    IoInMux I__1030 (
            .O(N__6737),
            .I(N__6734));
    LocalMux I__1029 (
            .O(N__6734),
            .I(N__6731));
    Span12Mux_s5_h I__1028 (
            .O(N__6731),
            .I(N__6728));
    Odrv12 I__1027 (
            .O(N__6728),
            .I(\FSM_TEST_inst_slow.current_state_RNIR2L81_0Z0Z_1 ));
    InMux I__1026 (
            .O(N__6725),
            .I(N__6722));
    LocalMux I__1025 (
            .O(N__6722),
            .I(\FSM_TEST_inst_slow.current_state_cnv_0_1 ));
    InMux I__1024 (
            .O(N__6719),
            .I(N__6709));
    InMux I__1023 (
            .O(N__6718),
            .I(N__6709));
    InMux I__1022 (
            .O(N__6717),
            .I(N__6709));
    CascadeMux I__1021 (
            .O(N__6716),
            .I(N__6706));
    LocalMux I__1020 (
            .O(N__6709),
            .I(N__6703));
    InMux I__1019 (
            .O(N__6706),
            .I(N__6700));
    Span4Mux_h I__1018 (
            .O(N__6703),
            .I(N__6697));
    LocalMux I__1017 (
            .O(N__6700),
            .I(\FSM_TEST_inst_slow.N_108_li ));
    Odrv4 I__1016 (
            .O(N__6697),
            .I(\FSM_TEST_inst_slow.N_108_li ));
    InMux I__1015 (
            .O(N__6692),
            .I(N__6689));
    LocalMux I__1014 (
            .O(N__6689),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_7 ));
    InMux I__1013 (
            .O(N__6686),
            .I(N__6683));
    LocalMux I__1012 (
            .O(N__6683),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_8 ));
    InMux I__1011 (
            .O(N__6680),
            .I(N__6677));
    LocalMux I__1010 (
            .O(N__6677),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_9 ));
    InMux I__1009 (
            .O(N__6674),
            .I(N__6671));
    LocalMux I__1008 (
            .O(N__6671),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_53 ));
    InMux I__1007 (
            .O(N__6668),
            .I(N__6665));
    LocalMux I__1006 (
            .O(N__6665),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_10 ));
    InMux I__1005 (
            .O(N__6662),
            .I(N__6659));
    LocalMux I__1004 (
            .O(N__6659),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_11 ));
    InMux I__1003 (
            .O(N__6656),
            .I(N__6653));
    LocalMux I__1002 (
            .O(N__6653),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_54 ));
    InMux I__1001 (
            .O(N__6650),
            .I(N__6647));
    LocalMux I__1000 (
            .O(N__6647),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_55 ));
    InMux I__999 (
            .O(N__6644),
            .I(N__6641));
    LocalMux I__998 (
            .O(N__6641),
            .I(N__6638));
    Odrv12 I__997 (
            .O(N__6638),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_50 ));
    InMux I__996 (
            .O(N__6635),
            .I(N__6632));
    LocalMux I__995 (
            .O(N__6632),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_51 ));
    InMux I__994 (
            .O(N__6629),
            .I(N__6626));
    LocalMux I__993 (
            .O(N__6626),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_5 ));
    InMux I__992 (
            .O(N__6623),
            .I(N__6620));
    LocalMux I__991 (
            .O(N__6620),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_23 ));
    CascadeMux I__990 (
            .O(N__6617),
            .I(N__6613));
    InMux I__989 (
            .O(N__6616),
            .I(N__6610));
    InMux I__988 (
            .O(N__6613),
            .I(N__6606));
    LocalMux I__987 (
            .O(N__6610),
            .I(N__6603));
    InMux I__986 (
            .O(N__6609),
            .I(N__6599));
    LocalMux I__985 (
            .O(N__6606),
            .I(N__6596));
    Span4Mux_v I__984 (
            .O(N__6603),
            .I(N__6593));
    InMux I__983 (
            .O(N__6602),
            .I(N__6590));
    LocalMux I__982 (
            .O(N__6599),
            .I(N__6587));
    Odrv12 I__981 (
            .O(N__6596),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__980 (
            .O(N__6593),
            .I(CONSTANT_ONE_NET));
    LocalMux I__979 (
            .O(N__6590),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__978 (
            .O(N__6587),
            .I(CONSTANT_ONE_NET));
    InMux I__977 (
            .O(N__6578),
            .I(N__6575));
    LocalMux I__976 (
            .O(N__6575),
            .I(N__6572));
    Odrv4 I__975 (
            .O(N__6572),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_86 ));
    InMux I__974 (
            .O(N__6569),
            .I(N__6566));
    LocalMux I__973 (
            .O(N__6566),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_84 ));
    InMux I__972 (
            .O(N__6563),
            .I(N__6560));
    LocalMux I__971 (
            .O(N__6560),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_85 ));
    InMux I__970 (
            .O(N__6557),
            .I(N__6554));
    LocalMux I__969 (
            .O(N__6554),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_82 ));
    InMux I__968 (
            .O(N__6551),
            .I(N__6548));
    LocalMux I__967 (
            .O(N__6548),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_83 ));
    InMux I__966 (
            .O(N__6545),
            .I(N__6542));
    LocalMux I__965 (
            .O(N__6542),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_12 ));
    InMux I__964 (
            .O(N__6539),
            .I(N__6536));
    LocalMux I__963 (
            .O(N__6536),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_52 ));
    CascadeMux I__962 (
            .O(N__6533),
            .I(\FSM_TEST_inst_RAPIDA.counter_idlelde_2_cascade_ ));
    CascadeMux I__961 (
            .O(N__6530),
            .I(N__6525));
    CascadeMux I__960 (
            .O(N__6529),
            .I(N__6522));
    CascadeMux I__959 (
            .O(N__6528),
            .I(N__6517));
    InMux I__958 (
            .O(N__6525),
            .I(N__6510));
    InMux I__957 (
            .O(N__6522),
            .I(N__6510));
    InMux I__956 (
            .O(N__6521),
            .I(N__6510));
    InMux I__955 (
            .O(N__6520),
            .I(N__6507));
    InMux I__954 (
            .O(N__6517),
            .I(N__6504));
    LocalMux I__953 (
            .O(N__6510),
            .I(N__6501));
    LocalMux I__952 (
            .O(N__6507),
            .I(N__6498));
    LocalMux I__951 (
            .O(N__6504),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1 ));
    Odrv4 I__950 (
            .O(N__6501),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1 ));
    Odrv4 I__949 (
            .O(N__6498),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1 ));
    CascadeMux I__948 (
            .O(N__6491),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1_cascade_ ));
    InMux I__947 (
            .O(N__6488),
            .I(N__6475));
    InMux I__946 (
            .O(N__6487),
            .I(N__6475));
    InMux I__945 (
            .O(N__6486),
            .I(N__6475));
    InMux I__944 (
            .O(N__6485),
            .I(N__6475));
    InMux I__943 (
            .O(N__6484),
            .I(N__6472));
    LocalMux I__942 (
            .O(N__6475),
            .I(N__6467));
    LocalMux I__941 (
            .O(N__6472),
            .I(N__6467));
    Span4Mux_h I__940 (
            .O(N__6467),
            .I(N__6464));
    Odrv4 I__939 (
            .O(N__6464),
            .I(\FSM_TEST_inst_RAPIDA.N_126_1_i ));
    InMux I__938 (
            .O(N__6461),
            .I(N__6456));
    InMux I__937 (
            .O(N__6460),
            .I(N__6453));
    InMux I__936 (
            .O(N__6459),
            .I(N__6450));
    LocalMux I__935 (
            .O(N__6456),
            .I(N__6445));
    LocalMux I__934 (
            .O(N__6453),
            .I(N__6445));
    LocalMux I__933 (
            .O(N__6450),
            .I(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_1 ));
    Odrv4 I__932 (
            .O(N__6445),
            .I(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_1 ));
    CascadeMux I__931 (
            .O(N__6440),
            .I(N__6435));
    InMux I__930 (
            .O(N__6439),
            .I(N__6431));
    InMux I__929 (
            .O(N__6438),
            .I(N__6424));
    InMux I__928 (
            .O(N__6435),
            .I(N__6424));
    InMux I__927 (
            .O(N__6434),
            .I(N__6424));
    LocalMux I__926 (
            .O(N__6431),
            .I(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_2 ));
    LocalMux I__925 (
            .O(N__6424),
            .I(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_2 ));
    InMux I__924 (
            .O(N__6419),
            .I(N__6412));
    InMux I__923 (
            .O(N__6418),
            .I(N__6412));
    InMux I__922 (
            .O(N__6417),
            .I(N__6409));
    LocalMux I__921 (
            .O(N__6412),
            .I(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_0 ));
    LocalMux I__920 (
            .O(N__6409),
            .I(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_0 ));
    InMux I__919 (
            .O(N__6404),
            .I(N__6401));
    LocalMux I__918 (
            .O(N__6401),
            .I(\FSM_TEST_inst_RAPIDA.G_24_0_a4_1_5 ));
    InMux I__917 (
            .O(N__6398),
            .I(N__6395));
    LocalMux I__916 (
            .O(N__6395),
            .I(N__6392));
    Odrv4 I__915 (
            .O(N__6392),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_6 ));
    InMux I__914 (
            .O(N__6389),
            .I(N__6386));
    LocalMux I__913 (
            .O(N__6386),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_19 ));
    InMux I__912 (
            .O(N__6383),
            .I(N__6380));
    LocalMux I__911 (
            .O(N__6380),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_20 ));
    InMux I__910 (
            .O(N__6377),
            .I(N__6374));
    LocalMux I__909 (
            .O(N__6374),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_21 ));
    InMux I__908 (
            .O(N__6371),
            .I(N__6368));
    LocalMux I__907 (
            .O(N__6368),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_22 ));
    InMux I__906 (
            .O(N__6365),
            .I(N__6362));
    LocalMux I__905 (
            .O(N__6362),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_3 ));
    InMux I__904 (
            .O(N__6359),
            .I(N__6356));
    LocalMux I__903 (
            .O(N__6356),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_4 ));
    InMux I__902 (
            .O(N__6353),
            .I(N__6350));
    LocalMux I__901 (
            .O(N__6350),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_5 ));
    InMux I__900 (
            .O(N__6347),
            .I(N__6344));
    LocalMux I__899 (
            .O(N__6344),
            .I(\FSM_TEST_inst_RAPIDA.counter_idle_cry_3_THRU_CO ));
    InMux I__898 (
            .O(N__6341),
            .I(N__6338));
    LocalMux I__897 (
            .O(N__6338),
            .I(\FSM_TEST_inst_RAPIDA.flag_input_regZ0 ));
    InMux I__896 (
            .O(N__6335),
            .I(N__6332));
    LocalMux I__895 (
            .O(N__6332),
            .I(\FSM_TEST_inst_RAPIDA.G_24_0_a4_1_4 ));
    InMux I__894 (
            .O(N__6329),
            .I(N__6326));
    LocalMux I__893 (
            .O(N__6326),
            .I(\FSM_TEST_inst_RAPIDA.counter_idle_cry_1_THRU_CO ));
    InMux I__892 (
            .O(N__6323),
            .I(N__6320));
    LocalMux I__891 (
            .O(N__6320),
            .I(\FSM_TEST_inst_RAPIDA.counter_idle_cry_2_THRU_CO ));
    InMux I__890 (
            .O(N__6317),
            .I(N__6311));
    InMux I__889 (
            .O(N__6316),
            .I(N__6304));
    InMux I__888 (
            .O(N__6315),
            .I(N__6304));
    InMux I__887 (
            .O(N__6314),
            .I(N__6304));
    LocalMux I__886 (
            .O(N__6311),
            .I(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_4 ));
    LocalMux I__885 (
            .O(N__6304),
            .I(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_4 ));
    CascadeMux I__884 (
            .O(N__6299),
            .I(N__6295));
    InMux I__883 (
            .O(N__6298),
            .I(N__6290));
    InMux I__882 (
            .O(N__6295),
            .I(N__6283));
    InMux I__881 (
            .O(N__6294),
            .I(N__6283));
    InMux I__880 (
            .O(N__6293),
            .I(N__6283));
    LocalMux I__879 (
            .O(N__6290),
            .I(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_3 ));
    LocalMux I__878 (
            .O(N__6283),
            .I(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_3 ));
    CascadeMux I__877 (
            .O(N__6278),
            .I(N__6273));
    CascadeMux I__876 (
            .O(N__6277),
            .I(N__6270));
    InMux I__875 (
            .O(N__6276),
            .I(N__6267));
    InMux I__874 (
            .O(N__6273),
            .I(N__6264));
    InMux I__873 (
            .O(N__6270),
            .I(N__6261));
    LocalMux I__872 (
            .O(N__6267),
            .I(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_5 ));
    LocalMux I__871 (
            .O(N__6264),
            .I(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_5 ));
    LocalMux I__870 (
            .O(N__6261),
            .I(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_5 ));
    InMux I__869 (
            .O(N__6254),
            .I(N__6251));
    LocalMux I__868 (
            .O(N__6251),
            .I(N__6245));
    CascadeMux I__867 (
            .O(N__6250),
            .I(N__6241));
    CascadeMux I__866 (
            .O(N__6249),
            .I(N__6238));
    CascadeMux I__865 (
            .O(N__6248),
            .I(N__6234));
    Span4Mux_h I__864 (
            .O(N__6245),
            .I(N__6230));
    InMux I__863 (
            .O(N__6244),
            .I(N__6217));
    InMux I__862 (
            .O(N__6241),
            .I(N__6217));
    InMux I__861 (
            .O(N__6238),
            .I(N__6217));
    InMux I__860 (
            .O(N__6237),
            .I(N__6217));
    InMux I__859 (
            .O(N__6234),
            .I(N__6217));
    InMux I__858 (
            .O(N__6233),
            .I(N__6217));
    Odrv4 I__857 (
            .O(N__6230),
            .I(\FSM_TEST_inst_RAPIDA.current_state_d_i_2 ));
    LocalMux I__856 (
            .O(N__6217),
            .I(\FSM_TEST_inst_RAPIDA.current_state_d_i_2 ));
    InMux I__855 (
            .O(N__6212),
            .I(N__6207));
    InMux I__854 (
            .O(N__6211),
            .I(N__6204));
    InMux I__853 (
            .O(N__6210),
            .I(N__6201));
    LocalMux I__852 (
            .O(N__6207),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_7 ));
    LocalMux I__851 (
            .O(N__6204),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_7 ));
    LocalMux I__850 (
            .O(N__6201),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_7 ));
    CascadeMux I__849 (
            .O(N__6194),
            .I(N__6191));
    InMux I__848 (
            .O(N__6191),
            .I(N__6188));
    LocalMux I__847 (
            .O(N__6188),
            .I(\FSM_TEST_inst_slow.flag_input_regZ0 ));
    CascadeMux I__846 (
            .O(N__6185),
            .I(N__6181));
    InMux I__845 (
            .O(N__6184),
            .I(N__6177));
    InMux I__844 (
            .O(N__6181),
            .I(N__6174));
    InMux I__843 (
            .O(N__6180),
            .I(N__6171));
    LocalMux I__842 (
            .O(N__6177),
            .I(N__6168));
    LocalMux I__841 (
            .O(N__6174),
            .I(N__6165));
    LocalMux I__840 (
            .O(N__6171),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_6 ));
    Odrv4 I__839 (
            .O(N__6168),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_6 ));
    Odrv4 I__838 (
            .O(N__6165),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_6 ));
    InMux I__837 (
            .O(N__6158),
            .I(N__6155));
    LocalMux I__836 (
            .O(N__6155),
            .I(\FSM_TEST_inst_slow.current_state_RNO_3Z0Z_0 ));
    CascadeMux I__835 (
            .O(N__6152),
            .I(\FSM_TEST_inst_slow.current_state_RNO_4Z0Z_0_cascade_ ));
    InMux I__834 (
            .O(N__6149),
            .I(N__6146));
    LocalMux I__833 (
            .O(N__6146),
            .I(\FSM_TEST_inst_slow.current_state_RNO_5Z0Z_0 ));
    InMux I__832 (
            .O(N__6143),
            .I(N__6140));
    LocalMux I__831 (
            .O(N__6140),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_0 ));
    InMux I__830 (
            .O(N__6137),
            .I(N__6134));
    LocalMux I__829 (
            .O(N__6134),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_1 ));
    InMux I__828 (
            .O(N__6131),
            .I(N__6128));
    LocalMux I__827 (
            .O(N__6128),
            .I(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_2 ));
    InMux I__826 (
            .O(N__6125),
            .I(N__6118));
    InMux I__825 (
            .O(N__6124),
            .I(N__6118));
    InMux I__824 (
            .O(N__6123),
            .I(N__6115));
    LocalMux I__823 (
            .O(N__6118),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_0 ));
    LocalMux I__822 (
            .O(N__6115),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_0 ));
    InMux I__821 (
            .O(N__6110),
            .I(N__6107));
    LocalMux I__820 (
            .O(N__6107),
            .I(\FSM_TEST_inst_slow.counter_stat_cry_1_THRU_CO ));
    InMux I__819 (
            .O(N__6104),
            .I(N__6097));
    InMux I__818 (
            .O(N__6103),
            .I(N__6097));
    InMux I__817 (
            .O(N__6102),
            .I(N__6094));
    LocalMux I__816 (
            .O(N__6097),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_2 ));
    LocalMux I__815 (
            .O(N__6094),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_2 ));
    CascadeMux I__814 (
            .O(N__6089),
            .I(N__6086));
    InMux I__813 (
            .O(N__6086),
            .I(N__6083));
    LocalMux I__812 (
            .O(N__6083),
            .I(\FSM_TEST_inst_slow.counter_stat_cry_2_THRU_CO ));
    InMux I__811 (
            .O(N__6080),
            .I(N__6074));
    InMux I__810 (
            .O(N__6079),
            .I(N__6069));
    InMux I__809 (
            .O(N__6078),
            .I(N__6069));
    InMux I__808 (
            .O(N__6077),
            .I(N__6066));
    LocalMux I__807 (
            .O(N__6074),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_3 ));
    LocalMux I__806 (
            .O(N__6069),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_3 ));
    LocalMux I__805 (
            .O(N__6066),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_3 ));
    InMux I__804 (
            .O(N__6059),
            .I(N__6056));
    LocalMux I__803 (
            .O(N__6056),
            .I(\FSM_TEST_inst_slow.counter_stat_cry_0_THRU_CO ));
    InMux I__802 (
            .O(N__6053),
            .I(N__6048));
    InMux I__801 (
            .O(N__6052),
            .I(N__6045));
    InMux I__800 (
            .O(N__6051),
            .I(N__6042));
    LocalMux I__799 (
            .O(N__6048),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_1 ));
    LocalMux I__798 (
            .O(N__6045),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_1 ));
    LocalMux I__797 (
            .O(N__6042),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_1 ));
    InMux I__796 (
            .O(N__6035),
            .I(N__6032));
    LocalMux I__795 (
            .O(N__6032),
            .I(\FSM_TEST_inst_slow.counter_stat_cry_3_THRU_CO ));
    InMux I__794 (
            .O(N__6029),
            .I(N__6023));
    InMux I__793 (
            .O(N__6028),
            .I(N__6020));
    InMux I__792 (
            .O(N__6027),
            .I(N__6015));
    InMux I__791 (
            .O(N__6026),
            .I(N__6015));
    LocalMux I__790 (
            .O(N__6023),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_4 ));
    LocalMux I__789 (
            .O(N__6020),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_4 ));
    LocalMux I__788 (
            .O(N__6015),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_4 ));
    InMux I__787 (
            .O(N__6008),
            .I(N__6002));
    InMux I__786 (
            .O(N__6007),
            .I(N__5999));
    InMux I__785 (
            .O(N__6006),
            .I(N__5994));
    InMux I__784 (
            .O(N__6005),
            .I(N__5994));
    LocalMux I__783 (
            .O(N__6002),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_4 ));
    LocalMux I__782 (
            .O(N__5999),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_4 ));
    LocalMux I__781 (
            .O(N__5994),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_4 ));
    InMux I__780 (
            .O(N__5987),
            .I(N__5981));
    InMux I__779 (
            .O(N__5986),
            .I(N__5978));
    InMux I__778 (
            .O(N__5985),
            .I(N__5975));
    InMux I__777 (
            .O(N__5984),
            .I(N__5972));
    LocalMux I__776 (
            .O(N__5981),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_5 ));
    LocalMux I__775 (
            .O(N__5978),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_5 ));
    LocalMux I__774 (
            .O(N__5975),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_5 ));
    LocalMux I__773 (
            .O(N__5972),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_5 ));
    InMux I__772 (
            .O(N__5963),
            .I(N__5959));
    InMux I__771 (
            .O(N__5962),
            .I(N__5955));
    LocalMux I__770 (
            .O(N__5959),
            .I(N__5952));
    InMux I__769 (
            .O(N__5958),
            .I(N__5949));
    LocalMux I__768 (
            .O(N__5955),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_1 ));
    Odrv4 I__767 (
            .O(N__5952),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_1 ));
    LocalMux I__766 (
            .O(N__5949),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_1 ));
    InMux I__765 (
            .O(N__5942),
            .I(N__5939));
    LocalMux I__764 (
            .O(N__5939),
            .I(N__5936));
    Odrv4 I__763 (
            .O(N__5936),
            .I(\FSM_TEST_inst_RAPIDA.counter_idle_cry_0_THRU_CO ));
    CascadeMux I__762 (
            .O(N__5933),
            .I(\FSM_TEST_inst_RAPIDA.N_126_1_i_cascade_ ));
    InMux I__761 (
            .O(N__5930),
            .I(\FSM_TEST_inst_slow.counter_stat_cry_0 ));
    InMux I__760 (
            .O(N__5927),
            .I(\FSM_TEST_inst_slow.counter_stat_cry_1 ));
    InMux I__759 (
            .O(N__5924),
            .I(\FSM_TEST_inst_slow.counter_stat_cry_2 ));
    InMux I__758 (
            .O(N__5921),
            .I(\FSM_TEST_inst_slow.counter_stat_cry_3 ));
    InMux I__757 (
            .O(N__5918),
            .I(\FSM_TEST_inst_slow.counter_stat_cry_4 ));
    InMux I__756 (
            .O(N__5915),
            .I(\FSM_TEST_inst_slow.counter_stat_cry_5 ));
    CascadeMux I__755 (
            .O(N__5912),
            .I(N__5907));
    CascadeMux I__754 (
            .O(N__5911),
            .I(N__5904));
    CascadeMux I__753 (
            .O(N__5910),
            .I(N__5901));
    InMux I__752 (
            .O(N__5907),
            .I(N__5898));
    InMux I__751 (
            .O(N__5904),
            .I(N__5895));
    InMux I__750 (
            .O(N__5901),
            .I(N__5892));
    LocalMux I__749 (
            .O(N__5898),
            .I(N__5889));
    LocalMux I__748 (
            .O(N__5895),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_6 ));
    LocalMux I__747 (
            .O(N__5892),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_6 ));
    Odrv4 I__746 (
            .O(N__5889),
            .I(\FSM_TEST_inst_slow.counter_statZ0Z_6 ));
    CascadeMux I__745 (
            .O(N__5882),
            .I(\FSM_TEST_inst_slow.current_state_ns_0_a3_1_4_0_cascade_ ));
    InMux I__744 (
            .O(N__5879),
            .I(N__5876));
    LocalMux I__743 (
            .O(N__5876),
            .I(\FSM_TEST_inst_slow.current_state_ns_0_a3_1_5_0 ));
    InMux I__742 (
            .O(N__5873),
            .I(N__5870));
    LocalMux I__741 (
            .O(N__5870),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_2 ));
    InMux I__740 (
            .O(N__5867),
            .I(N__5864));
    LocalMux I__739 (
            .O(N__5864),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_3 ));
    InMux I__738 (
            .O(N__5861),
            .I(N__5858));
    LocalMux I__737 (
            .O(N__5858),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_80 ));
    InMux I__736 (
            .O(N__5855),
            .I(N__5852));
    LocalMux I__735 (
            .O(N__5852),
            .I(N__5849));
    Odrv4 I__734 (
            .O(N__5849),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_42 ));
    InMux I__733 (
            .O(N__5846),
            .I(N__5843));
    LocalMux I__732 (
            .O(N__5843),
            .I(N__5840));
    Odrv12 I__731 (
            .O(N__5840),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_70 ));
    InMux I__730 (
            .O(N__5837),
            .I(N__5834));
    LocalMux I__729 (
            .O(N__5834),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_45 ));
    InMux I__728 (
            .O(N__5831),
            .I(N__5828));
    LocalMux I__727 (
            .O(N__5828),
            .I(N__5825));
    Odrv4 I__726 (
            .O(N__5825),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_76 ));
    InMux I__725 (
            .O(N__5822),
            .I(N__5819));
    LocalMux I__724 (
            .O(N__5819),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_77 ));
    InMux I__723 (
            .O(N__5816),
            .I(N__5813));
    LocalMux I__722 (
            .O(N__5813),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_43 ));
    InMux I__721 (
            .O(N__5810),
            .I(N__5807));
    LocalMux I__720 (
            .O(N__5807),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_44 ));
    InMux I__719 (
            .O(N__5804),
            .I(N__5801));
    LocalMux I__718 (
            .O(N__5801),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_78 ));
    InMux I__717 (
            .O(N__5798),
            .I(N__5795));
    LocalMux I__716 (
            .O(N__5795),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_79 ));
    InMux I__715 (
            .O(N__5792),
            .I(N__5789));
    LocalMux I__714 (
            .O(N__5789),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_13 ));
    InMux I__713 (
            .O(N__5786),
            .I(N__5783));
    LocalMux I__712 (
            .O(N__5783),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_0 ));
    InMux I__711 (
            .O(N__5780),
            .I(N__5777));
    LocalMux I__710 (
            .O(N__5777),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_81 ));
    InMux I__709 (
            .O(N__5774),
            .I(N__5771));
    LocalMux I__708 (
            .O(N__5771),
            .I(N__5768));
    Odrv4 I__707 (
            .O(N__5768),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_46 ));
    InMux I__706 (
            .O(N__5765),
            .I(N__5762));
    LocalMux I__705 (
            .O(N__5762),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_4 ));
    InMux I__704 (
            .O(N__5759),
            .I(N__5756));
    LocalMux I__703 (
            .O(N__5756),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_1 ));
    CascadeMux I__702 (
            .O(N__5753),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2Z0Z_1_cascade_ ));
    InMux I__701 (
            .O(N__5750),
            .I(N__5745));
    InMux I__700 (
            .O(N__5749),
            .I(N__5742));
    InMux I__699 (
            .O(N__5748),
            .I(N__5739));
    LocalMux I__698 (
            .O(N__5745),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_0 ));
    LocalMux I__697 (
            .O(N__5742),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_0 ));
    LocalMux I__696 (
            .O(N__5739),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_0 ));
    InMux I__695 (
            .O(N__5732),
            .I(N__5729));
    LocalMux I__694 (
            .O(N__5729),
            .I(\FSM_TEST_inst_RAPIDA.counter_stat_cry_0_THRU_CO ));
    CascadeMux I__693 (
            .O(N__5726),
            .I(N__5721));
    InMux I__692 (
            .O(N__5725),
            .I(N__5715));
    InMux I__691 (
            .O(N__5724),
            .I(N__5704));
    InMux I__690 (
            .O(N__5721),
            .I(N__5704));
    InMux I__689 (
            .O(N__5720),
            .I(N__5704));
    InMux I__688 (
            .O(N__5719),
            .I(N__5704));
    InMux I__687 (
            .O(N__5718),
            .I(N__5704));
    LocalMux I__686 (
            .O(N__5715),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2Z0Z_1 ));
    LocalMux I__685 (
            .O(N__5704),
            .I(\FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2Z0Z_1 ));
    CascadeMux I__684 (
            .O(N__5699),
            .I(N__5696));
    InMux I__683 (
            .O(N__5696),
            .I(N__5693));
    LocalMux I__682 (
            .O(N__5693),
            .I(\FSM_TEST_inst_RAPIDA.counter_stat_cry_1_THRU_CO ));
    InMux I__681 (
            .O(N__5690),
            .I(N__5685));
    InMux I__680 (
            .O(N__5689),
            .I(N__5682));
    InMux I__679 (
            .O(N__5688),
            .I(N__5679));
    LocalMux I__678 (
            .O(N__5685),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_2 ));
    LocalMux I__677 (
            .O(N__5682),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_2 ));
    LocalMux I__676 (
            .O(N__5679),
            .I(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_2 ));
    InMux I__675 (
            .O(N__5672),
            .I(\FSM_TEST_inst_RAPIDA.counter_idle_cry_0 ));
    InMux I__674 (
            .O(N__5669),
            .I(\FSM_TEST_inst_RAPIDA.counter_idle_cry_1 ));
    InMux I__673 (
            .O(N__5666),
            .I(\FSM_TEST_inst_RAPIDA.counter_idle_cry_2 ));
    InMux I__672 (
            .O(N__5663),
            .I(\FSM_TEST_inst_RAPIDA.counter_idle_cry_3 ));
    InMux I__671 (
            .O(N__5660),
            .I(\FSM_TEST_inst_RAPIDA.counter_idle_cry_4 ));
    InMux I__670 (
            .O(N__5657),
            .I(N__5645));
    InMux I__669 (
            .O(N__5656),
            .I(N__5645));
    InMux I__668 (
            .O(N__5655),
            .I(N__5645));
    InMux I__667 (
            .O(N__5654),
            .I(N__5645));
    LocalMux I__666 (
            .O(N__5645),
            .I(N__5638));
    InMux I__665 (
            .O(N__5644),
            .I(N__5629));
    InMux I__664 (
            .O(N__5643),
            .I(N__5629));
    InMux I__663 (
            .O(N__5642),
            .I(N__5629));
    InMux I__662 (
            .O(N__5641),
            .I(N__5629));
    Odrv4 I__661 (
            .O(N__5638),
            .I(\FSM_TEST_inst_slow.N_134_1_i ));
    LocalMux I__660 (
            .O(N__5629),
            .I(\FSM_TEST_inst_slow.N_134_1_i ));
    InMux I__659 (
            .O(N__5624),
            .I(N__5619));
    InMux I__658 (
            .O(N__5623),
            .I(N__5616));
    InMux I__657 (
            .O(N__5622),
            .I(N__5613));
    LocalMux I__656 (
            .O(N__5619),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_4 ));
    LocalMux I__655 (
            .O(N__5616),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_4 ));
    LocalMux I__654 (
            .O(N__5613),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_4 ));
    InMux I__653 (
            .O(N__5606),
            .I(N__5601));
    InMux I__652 (
            .O(N__5605),
            .I(N__5598));
    InMux I__651 (
            .O(N__5604),
            .I(N__5595));
    LocalMux I__650 (
            .O(N__5601),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_3 ));
    LocalMux I__649 (
            .O(N__5598),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_3 ));
    LocalMux I__648 (
            .O(N__5595),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_3 ));
    InMux I__647 (
            .O(N__5588),
            .I(N__5585));
    LocalMux I__646 (
            .O(N__5585),
            .I(\FSM_TEST_inst_RAPIDA.counter_stat_cry_3_THRU_CO ));
    InMux I__645 (
            .O(N__5582),
            .I(N__5579));
    LocalMux I__644 (
            .O(N__5579),
            .I(\FSM_TEST_inst_RAPIDA.counter_stat_cry_4_THRU_CO ));
    InMux I__643 (
            .O(N__5576),
            .I(N__5573));
    LocalMux I__642 (
            .O(N__5573),
            .I(\FSM_TEST_inst_RAPIDA.counter_stat_cry_2_THRU_CO ));
    CascadeMux I__641 (
            .O(N__5570),
            .I(\FSM_TEST_inst_RAPIDA.counter_statlde_0_cascade_ ));
    InMux I__640 (
            .O(N__5567),
            .I(\FSM_TEST_inst_slow.counter_idle_cry_1 ));
    InMux I__639 (
            .O(N__5564),
            .I(\FSM_TEST_inst_slow.counter_idle_cry_2 ));
    InMux I__638 (
            .O(N__5561),
            .I(\FSM_TEST_inst_slow.counter_idle_cry_3 ));
    InMux I__637 (
            .O(N__5558),
            .I(\FSM_TEST_inst_slow.counter_idle_cry_4 ));
    InMux I__636 (
            .O(N__5555),
            .I(\FSM_TEST_inst_slow.counter_idle_cry_5 ));
    InMux I__635 (
            .O(N__5552),
            .I(\FSM_TEST_inst_slow.counter_idle_cry_6 ));
    CEMux I__634 (
            .O(N__5549),
            .I(N__5546));
    LocalMux I__633 (
            .O(N__5546),
            .I(N__5543));
    Span4Mux_h I__632 (
            .O(N__5543),
            .I(N__5540));
    Odrv4 I__631 (
            .O(N__5540),
            .I(\FSM_TEST_inst_slow.counter_idle_RNIHR3A2Z0Z_7 ));
    InMux I__630 (
            .O(N__5537),
            .I(N__5533));
    InMux I__629 (
            .O(N__5536),
            .I(N__5530));
    LocalMux I__628 (
            .O(N__5533),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_1 ));
    LocalMux I__627 (
            .O(N__5530),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_1 ));
    InMux I__626 (
            .O(N__5525),
            .I(N__5521));
    InMux I__625 (
            .O(N__5524),
            .I(N__5518));
    LocalMux I__624 (
            .O(N__5521),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_2 ));
    LocalMux I__623 (
            .O(N__5518),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_2 ));
    CascadeMux I__622 (
            .O(N__5513),
            .I(N__5510));
    InMux I__621 (
            .O(N__5510),
            .I(N__5506));
    InMux I__620 (
            .O(N__5509),
            .I(N__5502));
    LocalMux I__619 (
            .O(N__5506),
            .I(N__5499));
    InMux I__618 (
            .O(N__5505),
            .I(N__5496));
    LocalMux I__617 (
            .O(N__5502),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_5 ));
    Odrv4 I__616 (
            .O(N__5499),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_5 ));
    LocalMux I__615 (
            .O(N__5496),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_5 ));
    InMux I__614 (
            .O(N__5489),
            .I(N__5485));
    InMux I__613 (
            .O(N__5488),
            .I(N__5482));
    LocalMux I__612 (
            .O(N__5485),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_0 ));
    LocalMux I__611 (
            .O(N__5482),
            .I(\FSM_TEST_inst_slow.counter_idleZ0Z_0 ));
    InMux I__610 (
            .O(N__5477),
            .I(N__5474));
    LocalMux I__609 (
            .O(N__5474),
            .I(\FSM_TEST_inst_slow.N_109_0 ));
    CascadeMux I__608 (
            .O(N__5471),
            .I(N__5468));
    InMux I__607 (
            .O(N__5468),
            .I(N__5460));
    InMux I__606 (
            .O(N__5467),
            .I(N__5460));
    InMux I__605 (
            .O(N__5466),
            .I(N__5455));
    InMux I__604 (
            .O(N__5465),
            .I(N__5455));
    LocalMux I__603 (
            .O(N__5460),
            .I(\FSM_TEST_inst_slow.counter_dinZ0Z_0 ));
    LocalMux I__602 (
            .O(N__5455),
            .I(\FSM_TEST_inst_slow.counter_dinZ0Z_0 ));
    CascadeMux I__601 (
            .O(N__5450),
            .I(N__5446));
    InMux I__600 (
            .O(N__5449),
            .I(N__5442));
    InMux I__599 (
            .O(N__5446),
            .I(N__5437));
    InMux I__598 (
            .O(N__5445),
            .I(N__5437));
    LocalMux I__597 (
            .O(N__5442),
            .I(N__5432));
    LocalMux I__596 (
            .O(N__5437),
            .I(N__5432));
    Odrv4 I__595 (
            .O(N__5432),
            .I(\FSM_TEST_inst_slow.counter_dinZ1Z_1 ));
    CascadeMux I__594 (
            .O(N__5429),
            .I(\FSM_TEST_inst_slow.N_134_1_cascade_ ));
    InMux I__593 (
            .O(N__5426),
            .I(N__5423));
    LocalMux I__592 (
            .O(N__5423),
            .I(N__5420));
    Odrv4 I__591 (
            .O(N__5420),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_15 ));
    CascadeMux I__590 (
            .O(N__5417),
            .I(N__5414));
    InMux I__589 (
            .O(N__5414),
            .I(N__5411));
    LocalMux I__588 (
            .O(N__5411),
            .I(N__5408));
    Span4Mux_v I__587 (
            .O(N__5408),
            .I(N__5405));
    Odrv4 I__586 (
            .O(N__5405),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_87 ));
    InMux I__585 (
            .O(N__5402),
            .I(N__5399));
    LocalMux I__584 (
            .O(N__5399),
            .I(\FSM_TEST_inst_slow.G_31_1 ));
    CascadeMux I__583 (
            .O(N__5396),
            .I(\FSM_TEST_inst_slow.counter_statlde_0_cascade_ ));
    CEMux I__582 (
            .O(N__5393),
            .I(N__5390));
    LocalMux I__581 (
            .O(N__5390),
            .I(N__5386));
    CEMux I__580 (
            .O(N__5389),
            .I(N__5383));
    Span4Mux_h I__579 (
            .O(N__5386),
            .I(N__5380));
    LocalMux I__578 (
            .O(N__5383),
            .I(N__5377));
    Span4Mux_h I__577 (
            .O(N__5380),
            .I(N__5374));
    Odrv4 I__576 (
            .O(N__5377),
            .I(\FSM_TEST_inst_slow.current_state_RNIR2L81Z0Z_1 ));
    Odrv4 I__575 (
            .O(N__5374),
            .I(\FSM_TEST_inst_slow.current_state_RNIR2L81Z0Z_1 ));
    InMux I__574 (
            .O(N__5369),
            .I(bfn_10_18_0_));
    InMux I__573 (
            .O(N__5366),
            .I(\FSM_TEST_inst_slow.counter_idle_cry_0 ));
    InMux I__572 (
            .O(N__5363),
            .I(N__5360));
    LocalMux I__571 (
            .O(N__5360),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_26 ));
    InMux I__570 (
            .O(N__5357),
            .I(N__5354));
    LocalMux I__569 (
            .O(N__5354),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_29 ));
    InMux I__568 (
            .O(N__5351),
            .I(N__5348));
    LocalMux I__567 (
            .O(N__5348),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_23 ));
    InMux I__566 (
            .O(N__5345),
            .I(N__5342));
    LocalMux I__565 (
            .O(N__5342),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_24 ));
    InMux I__564 (
            .O(N__5339),
            .I(N__5336));
    LocalMux I__563 (
            .O(N__5336),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_27 ));
    InMux I__562 (
            .O(N__5333),
            .I(N__5330));
    LocalMux I__561 (
            .O(N__5330),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_28 ));
    InMux I__560 (
            .O(N__5327),
            .I(N__5324));
    LocalMux I__559 (
            .O(N__5324),
            .I(N__5321));
    Odrv4 I__558 (
            .O(N__5321),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_47 ));
    InMux I__557 (
            .O(N__5318),
            .I(N__5315));
    LocalMux I__556 (
            .O(N__5315),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_73 ));
    InMux I__555 (
            .O(N__5312),
            .I(N__5309));
    LocalMux I__554 (
            .O(N__5309),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_74 ));
    InMux I__553 (
            .O(N__5306),
            .I(N__5303));
    LocalMux I__552 (
            .O(N__5303),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_75 ));
    InMux I__551 (
            .O(N__5300),
            .I(N__5297));
    LocalMux I__550 (
            .O(N__5297),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_15 ));
    InMux I__549 (
            .O(N__5294),
            .I(N__5291));
    LocalMux I__548 (
            .O(N__5291),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_14 ));
    InMux I__547 (
            .O(N__5288),
            .I(N__5285));
    LocalMux I__546 (
            .O(N__5285),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_22 ));
    InMux I__545 (
            .O(N__5282),
            .I(N__5279));
    LocalMux I__544 (
            .O(N__5279),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_20 ));
    InMux I__543 (
            .O(N__5276),
            .I(N__5273));
    LocalMux I__542 (
            .O(N__5273),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_21 ));
    InMux I__541 (
            .O(N__5270),
            .I(N__5267));
    LocalMux I__540 (
            .O(N__5267),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_18 ));
    InMux I__539 (
            .O(N__5264),
            .I(N__5261));
    LocalMux I__538 (
            .O(N__5261),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_19 ));
    InMux I__537 (
            .O(N__5258),
            .I(N__5255));
    LocalMux I__536 (
            .O(N__5255),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_25 ));
    InMux I__535 (
            .O(N__5252),
            .I(N__5249));
    LocalMux I__534 (
            .O(N__5249),
            .I(\FSM_TEST_inst_slow.CLK_uC_6jZ0Z_0 ));
    InMux I__533 (
            .O(N__5246),
            .I(N__5243));
    LocalMux I__532 (
            .O(N__5243),
            .I(N__5240));
    Odrv4 I__531 (
            .O(N__5240),
            .I(\FSM_TEST_inst_slow.CLK_uC_6gZ0Z_0 ));
    InMux I__530 (
            .O(N__5237),
            .I(N__5234));
    LocalMux I__529 (
            .O(N__5234),
            .I(\FSM_TEST_inst_slow.CLK_uC_6hZ0Z_0 ));
    InMux I__528 (
            .O(N__5231),
            .I(\FSM_TEST_inst_RAPIDA.counter_stat_cry_0 ));
    InMux I__527 (
            .O(N__5228),
            .I(\FSM_TEST_inst_RAPIDA.counter_stat_cry_1 ));
    InMux I__526 (
            .O(N__5225),
            .I(\FSM_TEST_inst_RAPIDA.counter_stat_cry_2 ));
    InMux I__525 (
            .O(N__5222),
            .I(\FSM_TEST_inst_RAPIDA.counter_stat_cry_3 ));
    InMux I__524 (
            .O(N__5219),
            .I(\FSM_TEST_inst_RAPIDA.counter_stat_cry_4 ));
    InMux I__523 (
            .O(N__5216),
            .I(\FSM_TEST_inst_RAPIDA.counter_stat_cry_5 ));
    InMux I__522 (
            .O(N__5213),
            .I(N__5210));
    LocalMux I__521 (
            .O(N__5210),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_7 ));
    InMux I__520 (
            .O(N__5207),
            .I(N__5204));
    LocalMux I__519 (
            .O(N__5204),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_8 ));
    InMux I__518 (
            .O(N__5201),
            .I(N__5198));
    LocalMux I__517 (
            .O(N__5198),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_9 ));
    InMux I__516 (
            .O(N__5195),
            .I(N__5192));
    LocalMux I__515 (
            .O(N__5192),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_10 ));
    InMux I__514 (
            .O(N__5189),
            .I(N__5186));
    LocalMux I__513 (
            .O(N__5186),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_0 ));
    InMux I__512 (
            .O(N__5183),
            .I(N__5180));
    LocalMux I__511 (
            .O(N__5180),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_1 ));
    InMux I__510 (
            .O(N__5177),
            .I(N__5174));
    LocalMux I__509 (
            .O(N__5174),
            .I(\FSM_TEST_inst_slow.CLK_uC_6iZ0Z_0 ));
    InMux I__508 (
            .O(N__5171),
            .I(N__5168));
    LocalMux I__507 (
            .O(N__5168),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_13 ));
    InMux I__506 (
            .O(N__5165),
            .I(N__5162));
    LocalMux I__505 (
            .O(N__5162),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_3 ));
    InMux I__504 (
            .O(N__5159),
            .I(N__5156));
    LocalMux I__503 (
            .O(N__5156),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_2 ));
    InMux I__502 (
            .O(N__5153),
            .I(N__5150));
    LocalMux I__501 (
            .O(N__5150),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_11 ));
    InMux I__500 (
            .O(N__5147),
            .I(N__5144));
    LocalMux I__499 (
            .O(N__5144),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_14 ));
    InMux I__498 (
            .O(N__5141),
            .I(N__5138));
    LocalMux I__497 (
            .O(N__5138),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_4 ));
    InMux I__496 (
            .O(N__5135),
            .I(N__5132));
    LocalMux I__495 (
            .O(N__5132),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_5 ));
    InMux I__494 (
            .O(N__5129),
            .I(N__5126));
    LocalMux I__493 (
            .O(N__5126),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_6 ));
    InMux I__492 (
            .O(N__5123),
            .I(N__5120));
    LocalMux I__491 (
            .O(N__5120),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_30 ));
    InMux I__490 (
            .O(N__5117),
            .I(N__5114));
    LocalMux I__489 (
            .O(N__5114),
            .I(N__5111));
    Odrv4 I__488 (
            .O(N__5111),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_71 ));
    InMux I__487 (
            .O(N__5108),
            .I(N__5105));
    LocalMux I__486 (
            .O(N__5105),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_31 ));
    InMux I__485 (
            .O(N__5102),
            .I(N__5099));
    LocalMux I__484 (
            .O(N__5099),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_32 ));
    InMux I__483 (
            .O(N__5096),
            .I(N__5093));
    LocalMux I__482 (
            .O(N__5093),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_72 ));
    InMux I__481 (
            .O(N__5090),
            .I(N__5087));
    LocalMux I__480 (
            .O(N__5087),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_41 ));
    InMux I__479 (
            .O(N__5084),
            .I(N__5081));
    LocalMux I__478 (
            .O(N__5081),
            .I(N__5078));
    Span4Mux_v I__477 (
            .O(N__5078),
            .I(N__5075));
    Odrv4 I__476 (
            .O(N__5075),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_39 ));
    InMux I__475 (
            .O(N__5072),
            .I(N__5069));
    LocalMux I__474 (
            .O(N__5069),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_40 ));
    InMux I__473 (
            .O(N__5066),
            .I(N__5063));
    LocalMux I__472 (
            .O(N__5063),
            .I(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_12 ));
    InMux I__471 (
            .O(N__5060),
            .I(N__5057));
    LocalMux I__470 (
            .O(N__5057),
            .I(\FSM_TEST_inst_slow.CLK_uC_6eZ0Z_0 ));
    InMux I__469 (
            .O(N__5054),
            .I(N__5051));
    LocalMux I__468 (
            .O(N__5051),
            .I(\FSM_TEST_inst_slow.CLK_uC_6fZ0Z_0 ));
    InMux I__467 (
            .O(N__5048),
            .I(N__5045));
    LocalMux I__466 (
            .O(N__5045),
            .I(\FSM_TEST_inst_slow.CLK_uC_3_0_0 ));
    InMux I__465 (
            .O(N__5042),
            .I(N__5039));
    LocalMux I__464 (
            .O(N__5039),
            .I(\FSM_TEST_inst_slow.CLK_uC_4_0_0 ));
    InMux I__463 (
            .O(N__5036),
            .I(N__5033));
    LocalMux I__462 (
            .O(N__5033),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_16 ));
    InMux I__461 (
            .O(N__5030),
            .I(N__5027));
    LocalMux I__460 (
            .O(N__5027),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_17 ));
    InMux I__459 (
            .O(N__5024),
            .I(N__5021));
    LocalMux I__458 (
            .O(N__5021),
            .I(N__5018));
    Odrv4 I__457 (
            .O(N__5018),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_33 ));
    InMux I__456 (
            .O(N__5015),
            .I(N__5012));
    LocalMux I__455 (
            .O(N__5012),
            .I(N__5009));
    Odrv4 I__454 (
            .O(N__5009),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_48 ));
    CascadeMux I__453 (
            .O(N__5006),
            .I(N__5002));
    InMux I__452 (
            .O(N__5005),
            .I(N__4997));
    InMux I__451 (
            .O(N__5002),
            .I(N__4997));
    LocalMux I__450 (
            .O(N__4997),
            .I(\FSM_TEST_inst_slow.CLK_uCZ0 ));
    InMux I__449 (
            .O(N__4994),
            .I(N__4991));
    LocalMux I__448 (
            .O(N__4991),
            .I(\FSM_TEST_inst_slow.CLK_uC_6c_0_0 ));
    InMux I__447 (
            .O(N__4988),
            .I(N__4985));
    LocalMux I__446 (
            .O(N__4985),
            .I(\FSM_TEST_inst_slow.CLK_uC_6b_0_0 ));
    InMux I__445 (
            .O(N__4982),
            .I(N__4979));
    LocalMux I__444 (
            .O(N__4979),
            .I(\FSM_TEST_inst_slow.CLK_uC_2_0_0 ));
    InMux I__443 (
            .O(N__4976),
            .I(N__4973));
    LocalMux I__442 (
            .O(N__4973),
            .I(\FSM_TEST_inst_slow.CLK_uC_5_0_0 ));
    InMux I__441 (
            .O(N__4970),
            .I(N__4967));
    LocalMux I__440 (
            .O(N__4967),
            .I(\FSM_TEST_inst_slow.CLK_uC_6_0_0 ));
    InMux I__439 (
            .O(N__4964),
            .I(N__4961));
    LocalMux I__438 (
            .O(N__4961),
            .I(\FSM_TEST_inst_slow.CLK_uC_6dZ0Z_0 ));
    IoInMux I__437 (
            .O(N__4958),
            .I(N__4955));
    LocalMux I__436 (
            .O(N__4955),
            .I(N__4952));
    Span4Mux_s3_v I__435 (
            .O(N__4952),
            .I(N__4949));
    Span4Mux_h I__434 (
            .O(N__4949),
            .I(N__4946));
    Odrv4 I__433 (
            .O(N__4946),
            .I(DYNCNF_i_0));
    InMux I__432 (
            .O(N__4943),
            .I(N__4940));
    LocalMux I__431 (
            .O(N__4940),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_49 ));
    InMux I__430 (
            .O(N__4937),
            .I(N__4934));
    LocalMux I__429 (
            .O(N__4934),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_38 ));
    InMux I__428 (
            .O(N__4931),
            .I(N__4928));
    LocalMux I__427 (
            .O(N__4928),
            .I(N__4925));
    Odrv4 I__426 (
            .O(N__4925),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_34 ));
    InMux I__425 (
            .O(N__4922),
            .I(N__4919));
    LocalMux I__424 (
            .O(N__4919),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_35 ));
    InMux I__423 (
            .O(N__4916),
            .I(N__4913));
    LocalMux I__422 (
            .O(N__4913),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_36 ));
    InMux I__421 (
            .O(N__4910),
            .I(N__4907));
    LocalMux I__420 (
            .O(N__4907),
            .I(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_37 ));
    IoInMux I__419 (
            .O(N__4904),
            .I(N__4901));
    LocalMux I__418 (
            .O(N__4901),
            .I(N__4898));
    IoSpan4Mux I__417 (
            .O(N__4898),
            .I(N__4895));
    Span4Mux_s3_v I__416 (
            .O(N__4895),
            .I(N__4892));
    Sp12to4 I__415 (
            .O(N__4892),
            .I(N__4889));
    Span12Mux_v I__414 (
            .O(N__4889),
            .I(N__4886));
    Span12Mux_v I__413 (
            .O(N__4886),
            .I(N__4883));
    Odrv12 I__412 (
            .O(N__4883),
            .I(CLK_c));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_18_0_));
    ICE_GB RST_N_ibuf_RNIBJGC_0 (
            .USERSIGNALTOGLOBALBUFFER(N__12008),
            .GLOBALBUFFEROUTPUT(RST_N_c_i_g));
    ICE_GB \FSM_TEST_inst_slow.current_state_RNIR2L81_1_1  (
            .USERSIGNALTOGLOBALBUFFER(N__6737),
            .GLOBALBUFFEROUTPUT(\FSM_TEST_inst_slow.N_374_g ));
    ICE_GB \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIKIU51_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__11885),
            .GLOBALBUFFEROUTPUT(\FSM_TEST_inst_RAPIDA.N_256_g ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_36_LC_6_17_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_36_LC_6_17_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_36_LC_6_17_3 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_36_LC_6_17_3  (
            .in0(N__7812),
            .in1(N__4922),
            .in2(_gnd_net_),
            .in3(N__8954),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10885),
            .ce(N__7310),
            .sr(N__10668));
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNIP1121_0_0_LC_7_1_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNIP1121_0_0_LC_7_1_2 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNIP1121_0_0_LC_7_1_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \config_register_latched_dec_inst.DYNCNF_1_RNIP1121_0_0_LC_7_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6791),
            .lcout(DYNCNF_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_50_LC_7_15_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_50_LC_7_15_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_50_LC_7_15_2 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_50_LC_7_15_2  (
            .in0(N__9049),
            .in1(_gnd_net_),
            .in2(N__7940),
            .in3(N__4943),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10868),
            .ce(N__7313),
            .sr(N__10671));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_49_LC_7_15_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_49_LC_7_15_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_49_LC_7_15_4 .LUT_INIT=16'b1111111110100101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_49_LC_7_15_4  (
            .in0(N__9048),
            .in1(_gnd_net_),
            .in2(N__7939),
            .in3(N__5015),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10868),
            .ce(N__7313),
            .sr(N__10671));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_34_LC_7_15_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_34_LC_7_15_7 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_34_LC_7_15_7 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_34_LC_7_15_7  (
            .in0(N__5024),
            .in1(N__7931),
            .in2(_gnd_net_),
            .in3(N__9047),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10868),
            .ce(N__7313),
            .sr(N__10671));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_71_LC_7_16_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_71_LC_7_16_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_71_LC_7_16_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_71_LC_7_16_5  (
            .in0(N__5846),
            .in1(N__7919),
            .in2(_gnd_net_),
            .in3(N__9046),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10874),
            .ce(N__7312),
            .sr(N__10669));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_39_LC_7_17_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_39_LC_7_17_0 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_39_LC_7_17_0 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_39_LC_7_17_0  (
            .in0(N__4937),
            .in1(N__7887),
            .in2(_gnd_net_),
            .in3(N__8953),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10880),
            .ce(N__7311),
            .sr(N__10664));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_38_LC_7_17_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_38_LC_7_17_1 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_38_LC_7_17_1 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_38_LC_7_17_1  (
            .in0(N__8952),
            .in1(N__4910),
            .in2(_gnd_net_),
            .in3(N__7888),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10880),
            .ce(N__7311),
            .sr(N__10664));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_35_LC_7_17_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_35_LC_7_17_2 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_35_LC_7_17_2 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_35_LC_7_17_2  (
            .in0(N__4931),
            .in1(N__7885),
            .in2(_gnd_net_),
            .in3(N__8950),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10880),
            .ce(N__7311),
            .sr(N__10664));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_37_LC_7_17_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_37_LC_7_17_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_37_LC_7_17_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_37_LC_7_17_6  (
            .in0(N__4916),
            .in1(N__7886),
            .in2(_gnd_net_),
            .in3(N__8951),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10880),
            .ce(N__7311),
            .sr(N__10664));
    defparam \FSM_TEST_inst_slow.CLK_uC_LC_7_18_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_LC_7_18_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_LC_7_18_0 .LUT_INIT=16'b1111011010010000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_LC_7_18_0  (
            .in0(N__7930),
            .in1(N__9045),
            .in2(N__5006),
            .in3(N__8546),
            .lcout(\FSM_TEST_inst_slow.CLK_uCZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10886),
            .ce(),
            .sr(N__10659));
    defparam \FSM_TEST_inst_slow.CLK_uC_6d_0_LC_7_18_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_6d_0_LC_7_18_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_6d_0_LC_7_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_6d_0_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4994),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_6dZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10886),
            .ce(),
            .sr(N__10659));
    defparam \FSM_TEST_inst_slow.CLK_uC_2_0_LC_7_18_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_2_0_LC_7_18_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_2_0_LC_7_18_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_2_0_LC_7_18_2  (
            .in0(N__5005),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10886),
            .ce(),
            .sr(N__10659));
    defparam \FSM_TEST_inst_slow.CLK_uC_6c_0_LC_7_18_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_6c_0_LC_7_18_3 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_6c_0_LC_7_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_6c_0_LC_7_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4988),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_6c_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10886),
            .ce(),
            .sr(N__10659));
    defparam \FSM_TEST_inst_slow.CLK_uC_5_0_LC_7_18_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_5_0_LC_7_18_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_5_0_LC_7_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_5_0_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5042),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10886),
            .ce(),
            .sr(N__10659));
    defparam \FSM_TEST_inst_slow.CLK_uC_6b_0_LC_7_18_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_6b_0_LC_7_18_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_6b_0_LC_7_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_6b_0_LC_7_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4970),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_6b_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10886),
            .ce(),
            .sr(N__10659));
    defparam \FSM_TEST_inst_slow.CLK_uC_3_0_LC_7_18_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_3_0_LC_7_18_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_3_0_LC_7_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_3_0_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4982),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10886),
            .ce(),
            .sr(N__10659));
    defparam \FSM_TEST_inst_slow.CLK_uC_6_0_LC_7_18_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_6_0_LC_7_18_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_6_0_LC_7_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_6_0_LC_7_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4976),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10886),
            .ce(),
            .sr(N__10659));
    defparam \FSM_TEST_inst_slow.CLK_uC_6e_0_LC_7_19_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_6e_0_LC_7_19_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_6e_0_LC_7_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_6e_0_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4964),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_6eZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10889),
            .ce(),
            .sr(N__10654));
    defparam \FSM_TEST_inst_slow.CLK_uC_6f_0_LC_7_19_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_6f_0_LC_7_19_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_6f_0_LC_7_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_6f_0_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5060),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_6fZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10889),
            .ce(),
            .sr(N__10654));
    defparam \FSM_TEST_inst_slow.CLK_uC_6g_0_LC_7_19_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_6g_0_LC_7_19_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_6g_0_LC_7_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_6g_0_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5054),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_6gZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10889),
            .ce(),
            .sr(N__10654));
    defparam \FSM_TEST_inst_slow.CLK_uC_4_0_LC_7_19_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_4_0_LC_7_19_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_4_0_LC_7_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_4_0_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5048),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10889),
            .ce(),
            .sr(N__10654));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_16_LC_9_13_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_16_LC_9_13_6 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_16_LC_9_13_6 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_16_LC_9_13_6  (
            .in0(N__5300),
            .in1(N__7909),
            .in2(_gnd_net_),
            .in3(N__9060),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10839),
            .ce(N__7323),
            .sr(N__10672));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_17_LC_9_13_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_17_LC_9_13_7 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_17_LC_9_13_7 .LUT_INIT=16'b1111111110100101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_17_LC_9_13_7  (
            .in0(N__9061),
            .in1(_gnd_net_),
            .in2(N__7938),
            .in3(N__5036),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10839),
            .ce(N__7323),
            .sr(N__10672));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_18_LC_9_14_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_18_LC_9_14_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_18_LC_9_14_0 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_18_LC_9_14_0  (
            .in0(N__9041),
            .in1(N__5030),
            .in2(_gnd_net_),
            .in3(N__7848),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10847),
            .ce(N__7319),
            .sr(N__10670));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_33_LC_9_15_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_33_LC_9_15_1 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_33_LC_9_15_1 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_33_LC_9_15_1  (
            .in0(N__5102),
            .in1(N__7841),
            .in2(_gnd_net_),
            .in3(N__9027),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10855),
            .ce(N__7316),
            .sr(N__10665));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_41_LC_9_15_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_41_LC_9_15_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_41_LC_9_15_2 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_41_LC_9_15_2  (
            .in0(N__9028),
            .in1(_gnd_net_),
            .in2(N__7921),
            .in3(N__5072),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10855),
            .ce(N__7316),
            .sr(N__10665));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_31_LC_9_15_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_31_LC_9_15_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_31_LC_9_15_4 .LUT_INIT=16'b1111111110100101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_31_LC_9_15_4  (
            .in0(N__9026),
            .in1(_gnd_net_),
            .in2(N__7920),
            .in3(N__5123),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10855),
            .ce(N__7316),
            .sr(N__10665));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_48_LC_9_15_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_48_LC_9_15_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_48_LC_9_15_6 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_48_LC_9_15_6  (
            .in0(N__9029),
            .in1(_gnd_net_),
            .in2(N__7922),
            .in3(N__5327),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10855),
            .ce(N__7316),
            .sr(N__10665));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_30_LC_9_15_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_30_LC_9_15_7 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_30_LC_9_15_7 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_30_LC_9_15_7  (
            .in0(N__5357),
            .in1(N__7837),
            .in2(_gnd_net_),
            .in3(N__9025),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10855),
            .ce(N__7316),
            .sr(N__10665));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_72_LC_9_16_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_72_LC_9_16_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_72_LC_9_16_0 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_72_LC_9_16_0  (
            .in0(N__8987),
            .in1(_gnd_net_),
            .in2(N__7917),
            .in3(N__5117),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10862),
            .ce(N__7314),
            .sr(N__10660));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_32_LC_9_16_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_32_LC_9_16_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_32_LC_9_16_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_32_LC_9_16_1  (
            .in0(N__5108),
            .in1(N__8984),
            .in2(_gnd_net_),
            .in3(N__7813),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10862),
            .ce(N__7314),
            .sr(N__10660));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_73_LC_9_16_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_73_LC_9_16_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_73_LC_9_16_2 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_73_LC_9_16_2  (
            .in0(N__8988),
            .in1(_gnd_net_),
            .in2(N__7918),
            .in3(N__5096),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10862),
            .ce(N__7314),
            .sr(N__10660));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_42_LC_9_16_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_42_LC_9_16_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_42_LC_9_16_4 .LUT_INIT=16'b1111111110100101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_42_LC_9_16_4  (
            .in0(N__8986),
            .in1(_gnd_net_),
            .in2(N__7916),
            .in3(N__5090),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10862),
            .ce(N__7314),
            .sr(N__10660));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_40_LC_9_16_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_40_LC_9_16_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_40_LC_9_16_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_40_LC_9_16_7  (
            .in0(N__5084),
            .in1(N__8985),
            .in2(_gnd_net_),
            .in3(N__7814),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10862),
            .ce(N__7314),
            .sr(N__10660));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_13_LC_9_17_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_13_LC_9_17_0 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_13_LC_9_17_0 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_13_LC_9_17_0  (
            .in0(N__7665),
            .in1(N__5066),
            .in2(_gnd_net_),
            .in3(N__8932),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10869),
            .ce(N__5393),
            .sr(N__10655));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_4_LC_9_17_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_4_LC_9_17_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_4_LC_9_17_1 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_4_LC_9_17_1  (
            .in0(N__8937),
            .in1(N__5165),
            .in2(_gnd_net_),
            .in3(N__7670),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10869),
            .ce(N__5393),
            .sr(N__10655));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_12_LC_9_17_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_12_LC_9_17_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_12_LC_9_17_2 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_12_LC_9_17_2  (
            .in0(N__7664),
            .in1(N__5153),
            .in2(_gnd_net_),
            .in3(N__8931),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10869),
            .ce(N__5393),
            .sr(N__10655));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_14_LC_9_17_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_14_LC_9_17_3 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_14_LC_9_17_3 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_14_LC_9_17_3  (
            .in0(N__8933),
            .in1(N__5171),
            .in2(_gnd_net_),
            .in3(N__7666),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10869),
            .ce(N__5393),
            .sr(N__10655));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_3_LC_9_17_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_3_LC_9_17_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_3_LC_9_17_4 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_3_LC_9_17_4  (
            .in0(N__7669),
            .in1(N__5159),
            .in2(_gnd_net_),
            .in3(N__8936),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10869),
            .ce(N__5393),
            .sr(N__10655));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_2_LC_9_17_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_2_LC_9_17_5 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_2_LC_9_17_5 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_2_LC_9_17_5  (
            .in0(N__8935),
            .in1(N__5183),
            .in2(_gnd_net_),
            .in3(N__7668),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10869),
            .ce(N__5393),
            .sr(N__10655));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_11_LC_9_17_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_11_LC_9_17_6 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_11_LC_9_17_6 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_11_LC_9_17_6  (
            .in0(N__7663),
            .in1(N__5195),
            .in2(_gnd_net_),
            .in3(N__8930),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10869),
            .ce(N__5393),
            .sr(N__10655));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_15_LC_9_17_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_15_LC_9_17_7 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_15_LC_9_17_7 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_15_LC_9_17_7  (
            .in0(N__8934),
            .in1(N__5147),
            .in2(_gnd_net_),
            .in3(N__7667),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10869),
            .ce(N__5393),
            .sr(N__10655));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_6_LC_9_18_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_6_LC_9_18_0 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_6_LC_9_18_0 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_6_LC_9_18_0  (
            .in0(N__9008),
            .in1(N__5135),
            .in2(_gnd_net_),
            .in3(N__7834),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10875),
            .ce(N__5389),
            .sr(N__10650));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_5_LC_9_18_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_5_LC_9_18_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_5_LC_9_18_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_5_LC_9_18_1  (
            .in0(N__5141),
            .in1(N__7831),
            .in2(_gnd_net_),
            .in3(N__9007),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10875),
            .ce(N__5389),
            .sr(N__10650));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_7_LC_9_18_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_7_LC_9_18_2 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_7_LC_9_18_2 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_7_LC_9_18_2  (
            .in0(N__9009),
            .in1(N__5129),
            .in2(_gnd_net_),
            .in3(N__7835),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10875),
            .ce(N__5389),
            .sr(N__10650));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_0_LC_9_18_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_0_LC_9_18_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_0_LC_9_18_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_0_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__7829),
            .in2(_gnd_net_),
            .in3(N__9004),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10875),
            .ce(N__5389),
            .sr(N__10650));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_8_LC_9_18_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_8_LC_9_18_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_8_LC_9_18_4 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_8_LC_9_18_4  (
            .in0(N__9010),
            .in1(N__5213),
            .in2(_gnd_net_),
            .in3(N__7836),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10875),
            .ce(N__5389),
            .sr(N__10650));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_9_LC_9_18_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_9_LC_9_18_5 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_9_LC_9_18_5 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_9_LC_9_18_5  (
            .in0(N__5207),
            .in1(N__7832),
            .in2(_gnd_net_),
            .in3(N__9011),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10875),
            .ce(N__5389),
            .sr(N__10650));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_10_LC_9_18_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_10_LC_9_18_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_10_LC_9_18_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_10_LC_9_18_6  (
            .in0(N__9005),
            .in1(N__5201),
            .in2(_gnd_net_),
            .in3(N__7833),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10875),
            .ce(N__5389),
            .sr(N__10650));
    defparam \FSM_TEST_inst_slow.bit_sequence_din_1_LC_9_18_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_1_LC_9_18_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_din_1_LC_9_18_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_din_1_LC_9_18_7  (
            .in0(N__5189),
            .in1(N__7830),
            .in2(_gnd_net_),
            .in3(N__9006),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_dinZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10875),
            .ce(N__5389),
            .sr(N__10650));
    defparam \FSM_TEST_inst_slow.counter_din_1_LC_9_19_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_din_1_LC_9_19_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_din_1_LC_9_19_0 .LUT_INIT=16'b0101110110000000;
    LogicCell40 \FSM_TEST_inst_slow.counter_din_1_LC_9_19_0  (
            .in0(N__7239),
            .in1(N__6718),
            .in2(N__5471),
            .in3(N__5449),
            .lcout(\FSM_TEST_inst_slow.counter_dinZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10881),
            .ce(),
            .sr(N__10646));
    defparam \FSM_TEST_inst_slow.counter_din_0_LC_9_19_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_din_0_LC_9_19_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_din_0_LC_9_19_1 .LUT_INIT=16'b0010001011001100;
    LogicCell40 \FSM_TEST_inst_slow.counter_din_0_LC_9_19_1  (
            .in0(N__6717),
            .in1(N__5467),
            .in2(_gnd_net_),
            .in3(N__7238),
            .lcout(\FSM_TEST_inst_slow.counter_dinZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10881),
            .ce(),
            .sr(N__10646));
    defparam \FSM_TEST_inst_slow.counter_din_3_LC_9_19_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_din_3_LC_9_19_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_din_3_LC_9_19_2 .LUT_INIT=16'b0101100011010000;
    LogicCell40 \FSM_TEST_inst_slow.counter_din_3_LC_9_19_2  (
            .in0(N__7240),
            .in1(N__6719),
            .in2(N__6942),
            .in3(N__5477),
            .lcout(\FSM_TEST_inst_slow.counter_dinZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10881),
            .ce(),
            .sr(N__10646));
    defparam \FSM_TEST_inst_slow.CLK_uC_6i_0_LC_9_19_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_6i_0_LC_9_19_3 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_6i_0_LC_9_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_6i_0_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5237),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_6iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10881),
            .ce(),
            .sr(N__10646));
    defparam \FSM_TEST_inst_slow.CLK_uC_6j_0_LC_9_19_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_6j_0_LC_9_19_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_6j_0_LC_9_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_6j_0_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5177),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_6jZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10881),
            .ce(),
            .sr(N__10646));
    defparam \FSM_TEST_inst_slow.CLK_uC_6k_0_LC_9_19_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_6k_0_LC_9_19_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_6k_0_LC_9_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_6k_0_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5252),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_6kZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10881),
            .ce(),
            .sr(N__10646));
    defparam \FSM_TEST_inst_slow.CLK_uC_6h_0_LC_9_19_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_6h_0_LC_9_19_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_6h_0_LC_9_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_6h_0_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5246),
            .lcout(\FSM_TEST_inst_slow.CLK_uC_6hZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10881),
            .ce(),
            .sr(N__10646));
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_c_0_LC_9_20_0 .C_ON=1'b1;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_c_0_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_c_0_LC_9_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_stat_cry_c_0_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__5748),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\FSM_TEST_inst_RAPIDA.counter_stat_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_0_THRU_LUT4_0_LC_9_20_1 .C_ON=1'b1;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_0_THRU_LUT4_0_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_0_THRU_LUT4_0_LC_9_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_stat_cry_0_THRU_LUT4_0_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__5958),
            .in2(_gnd_net_),
            .in3(N__5231),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_stat_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\FSM_TEST_inst_RAPIDA.counter_stat_cry_0 ),
            .carryout(\FSM_TEST_inst_RAPIDA.counter_stat_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_1_THRU_LUT4_0_LC_9_20_2 .C_ON=1'b1;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_1_THRU_LUT4_0_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_1_THRU_LUT4_0_LC_9_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_stat_cry_1_THRU_LUT4_0_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__5688),
            .in2(_gnd_net_),
            .in3(N__5228),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_stat_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\FSM_TEST_inst_RAPIDA.counter_stat_cry_1 ),
            .carryout(\FSM_TEST_inst_RAPIDA.counter_stat_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_2_THRU_LUT4_0_LC_9_20_3 .C_ON=1'b1;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_2_THRU_LUT4_0_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_2_THRU_LUT4_0_LC_9_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_stat_cry_2_THRU_LUT4_0_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__6985),
            .in2(_gnd_net_),
            .in3(N__5225),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_stat_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\FSM_TEST_inst_RAPIDA.counter_stat_cry_2 ),
            .carryout(\FSM_TEST_inst_RAPIDA.counter_stat_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_3_THRU_LUT4_0_LC_9_20_4 .C_ON=1'b1;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_3_THRU_LUT4_0_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_3_THRU_LUT4_0_LC_9_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_stat_cry_3_THRU_LUT4_0_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__6007),
            .in2(_gnd_net_),
            .in3(N__5222),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_stat_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\FSM_TEST_inst_RAPIDA.counter_stat_cry_3 ),
            .carryout(\FSM_TEST_inst_RAPIDA.counter_stat_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_4_THRU_LUT4_0_LC_9_20_5 .C_ON=1'b1;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_4_THRU_LUT4_0_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_cry_4_THRU_LUT4_0_LC_9_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_stat_cry_4_THRU_LUT4_0_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__5986),
            .in2(_gnd_net_),
            .in3(N__5219),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_stat_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\FSM_TEST_inst_RAPIDA.counter_stat_cry_4 ),
            .carryout(\FSM_TEST_inst_RAPIDA.counter_stat_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_6_LC_9_20_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_6_LC_9_20_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_6_LC_9_20_6 .LUT_INIT=16'b0011010001110000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_stat_6_LC_9_20_6  (
            .in0(N__6254),
            .in1(N__5725),
            .in2(N__7021),
            .in3(N__5216),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10887),
            .ce(),
            .sr(N__10641));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_87_LC_10_11_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_87_LC_10_11_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_87_LC_10_11_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_87_LC_10_11_4  (
            .in0(N__6578),
            .in1(N__7929),
            .in2(_gnd_net_),
            .in3(N__9062),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10821),
            .ce(N__7331),
            .sr(N__10673));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_15_LC_10_13_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_15_LC_10_13_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_15_LC_10_13_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_15_LC_10_13_1  (
            .in0(N__5294),
            .in1(N__7908),
            .in2(_gnd_net_),
            .in3(N__9051),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10826),
            .ce(N__7324),
            .sr(N__10666));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_14_LC_10_13_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_14_LC_10_13_7 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_14_LC_10_13_7 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_14_LC_10_13_7  (
            .in0(N__5792),
            .in1(N__7907),
            .in2(_gnd_net_),
            .in3(N__9050),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10826),
            .ce(N__7324),
            .sr(N__10666));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_23_LC_10_14_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_23_LC_10_14_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_23_LC_10_14_0 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_23_LC_10_14_0  (
            .in0(N__9024),
            .in1(N__5288),
            .in2(_gnd_net_),
            .in3(N__7881),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10832),
            .ce(N__7320),
            .sr(N__10661));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_20_LC_10_14_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_20_LC_10_14_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_20_LC_10_14_1 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_20_LC_10_14_1  (
            .in0(N__7878),
            .in1(N__5264),
            .in2(_gnd_net_),
            .in3(N__9021),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10832),
            .ce(N__7320),
            .sr(N__10661));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_22_LC_10_14_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_22_LC_10_14_3 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_22_LC_10_14_3 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_22_LC_10_14_3  (
            .in0(N__7880),
            .in1(N__5276),
            .in2(_gnd_net_),
            .in3(N__9023),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10832),
            .ce(N__7320),
            .sr(N__10661));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_21_LC_10_14_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_21_LC_10_14_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_21_LC_10_14_4 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_21_LC_10_14_4  (
            .in0(N__9022),
            .in1(N__5282),
            .in2(_gnd_net_),
            .in3(N__7879),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10832),
            .ce(N__7320),
            .sr(N__10661));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_19_LC_10_14_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_19_LC_10_14_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_19_LC_10_14_5 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_19_LC_10_14_5  (
            .in0(N__7877),
            .in1(N__5270),
            .in2(_gnd_net_),
            .in3(N__9020),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10832),
            .ce(N__7320),
            .sr(N__10661));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_26_LC_10_15_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_26_LC_10_15_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_26_LC_10_15_0 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_26_LC_10_15_0  (
            .in0(N__9015),
            .in1(_gnd_net_),
            .in2(N__7926),
            .in3(N__5258),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10841),
            .ce(N__7317),
            .sr(N__10656));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_25_LC_10_15_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_25_LC_10_15_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_25_LC_10_15_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_25_LC_10_15_1  (
            .in0(N__5345),
            .in1(N__7865),
            .in2(_gnd_net_),
            .in3(N__9014),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10841),
            .ce(N__7317),
            .sr(N__10656));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_27_LC_10_15_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_27_LC_10_15_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_27_LC_10_15_2 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_27_LC_10_15_2  (
            .in0(N__9016),
            .in1(_gnd_net_),
            .in2(N__7927),
            .in3(N__5363),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10841),
            .ce(N__7317),
            .sr(N__10656));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_29_LC_10_15_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_29_LC_10_15_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_29_LC_10_15_3 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_29_LC_10_15_3  (
            .in0(N__5333),
            .in1(N__7875),
            .in2(_gnd_net_),
            .in3(N__9018),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10841),
            .ce(N__7317),
            .sr(N__10656));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_24_LC_10_15_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_24_LC_10_15_5 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_24_LC_10_15_5 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_24_LC_10_15_5  (
            .in0(N__5351),
            .in1(N__7864),
            .in2(_gnd_net_),
            .in3(N__9013),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10841),
            .ce(N__7317),
            .sr(N__10656));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_28_LC_10_15_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_28_LC_10_15_6 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_28_LC_10_15_6 .LUT_INIT=16'b1111111110100101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_28_LC_10_15_6  (
            .in0(N__9017),
            .in1(_gnd_net_),
            .in2(N__7928),
            .in3(N__5339),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10841),
            .ce(N__7317),
            .sr(N__10656));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_47_LC_10_15_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_47_LC_10_15_7 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_47_LC_10_15_7 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_47_LC_10_15_7  (
            .in0(N__5774),
            .in1(N__7876),
            .in2(_gnd_net_),
            .in3(N__9019),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10841),
            .ce(N__7317),
            .sr(N__10656));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_76_LC_10_16_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_76_LC_10_16_0 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_76_LC_10_16_0 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_76_LC_10_16_0  (
            .in0(N__5306),
            .in1(N__7863),
            .in2(_gnd_net_),
            .in3(N__8983),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10849),
            .ce(N__7315),
            .sr(N__10651));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_74_LC_10_16_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_74_LC_10_16_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_74_LC_10_16_4 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_74_LC_10_16_4  (
            .in0(N__5318),
            .in1(N__7859),
            .in2(_gnd_net_),
            .in3(N__8981),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10849),
            .ce(N__7315),
            .sr(N__10651));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_75_LC_10_16_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_75_LC_10_16_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_75_LC_10_16_5 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_75_LC_10_16_5  (
            .in0(N__8982),
            .in1(_gnd_net_),
            .in2(N__7925),
            .in3(N__5312),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10849),
            .ce(N__7315),
            .sr(N__10651));
    defparam \FSM_TEST_inst_slow.current_state_RNIV6JP_2_1_LC_10_17_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNIV6JP_2_1_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNIV6JP_2_1_LC_10_17_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNIV6JP_2_1_LC_10_17_0  (
            .in0(N__7639),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8854),
            .lcout(),
            .ltout(\FSM_TEST_inst_slow.N_134_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.counter_idle_RNIHR3A2_7_LC_10_17_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_idle_RNIHR3A2_7_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.counter_idle_RNIHR3A2_7_LC_10_17_1 .LUT_INIT=16'b1101111100000000;
    LogicCell40 \FSM_TEST_inst_slow.counter_idle_RNIHR3A2_7_LC_10_17_1  (
            .in0(N__6211),
            .in1(N__5402),
            .in2(N__5429),
            .in3(N__7227),
            .lcout(\FSM_TEST_inst_slow.counter_idle_RNIHR3A2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.MOSI_er_LC_10_17_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.MOSI_er_LC_10_17_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.MOSI_er_LC_10_17_2 .LUT_INIT=16'b0100010010100000;
    LogicCell40 \FSM_TEST_inst_slow.MOSI_er_LC_10_17_2  (
            .in0(N__7644),
            .in1(N__5426),
            .in2(N__5417),
            .in3(N__8857),
            .lcout(mosi_slow),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10856),
            .ce(N__7241),
            .sr(N__10647));
    defparam \FSM_TEST_inst_slow.counter_idle_RNIMHOQ_3_LC_10_17_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_idle_RNIMHOQ_3_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.counter_idle_RNIMHOQ_3_LC_10_17_3 .LUT_INIT=16'b0000111100011111;
    LogicCell40 \FSM_TEST_inst_slow.counter_idle_RNIMHOQ_3_LC_10_17_3  (
            .in0(N__5605),
            .in1(N__5623),
            .in2(N__6185),
            .in3(N__5505),
            .lcout(\FSM_TEST_inst_slow.G_31_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.counter_stat_RNIE9EB1_6_LC_10_17_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_stat_RNIE9EB1_6_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.counter_stat_RNIE9EB1_6_LC_10_17_4 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \FSM_TEST_inst_slow.counter_stat_RNIE9EB1_6_LC_10_17_4  (
            .in0(N__9192),
            .in1(N__6026),
            .in2(N__5912),
            .in3(N__6077),
            .lcout(),
            .ltout(\FSM_TEST_inst_slow.counter_statlde_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.current_state_RNI9C3K2_1_LC_10_17_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNI9C3K2_1_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNI9C3K2_1_LC_10_17_5 .LUT_INIT=16'b1011111100000000;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNI9C3K2_1_LC_10_17_5  (
            .in0(N__8855),
            .in1(N__7640),
            .in2(N__5396),
            .in3(N__7225),
            .lcout(\FSM_TEST_inst_slow.current_state_RNI9C3K2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.current_state_RNIR2L81_1_LC_10_17_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNIR2L81_1_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNIR2L81_1_LC_10_17_6 .LUT_INIT=16'b1010101000001010;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNIR2L81_1_LC_10_17_6  (
            .in0(N__7226),
            .in1(_gnd_net_),
            .in2(N__7828),
            .in3(N__8856),
            .lcout(\FSM_TEST_inst_slow.current_state_RNIR2L81Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.current_state_RNO_7_0_LC_10_17_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNO_7_0_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNO_7_0_LC_10_17_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNO_7_0_LC_10_17_7  (
            .in0(N__6027),
            .in1(N__6052),
            .in2(N__9197),
            .in3(N__7638),
            .lcout(\FSM_TEST_inst_slow.current_state_ns_0_a3_1_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.counter_idle_0_LC_10_18_0 .C_ON=1'b1;
    defparam \FSM_TEST_inst_slow.counter_idle_0_LC_10_18_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_idle_0_LC_10_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \FSM_TEST_inst_slow.counter_idle_0_LC_10_18_0  (
            .in0(N__5654),
            .in1(N__5489),
            .in2(_gnd_net_),
            .in3(N__5369),
            .lcout(\FSM_TEST_inst_slow.counter_idleZ0Z_0 ),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\FSM_TEST_inst_slow.counter_idle_cry_0 ),
            .clk(N__10863),
            .ce(N__5549),
            .sr(N__10642));
    defparam \FSM_TEST_inst_slow.counter_idle_1_LC_10_18_1 .C_ON=1'b1;
    defparam \FSM_TEST_inst_slow.counter_idle_1_LC_10_18_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_idle_1_LC_10_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \FSM_TEST_inst_slow.counter_idle_1_LC_10_18_1  (
            .in0(N__5641),
            .in1(N__5537),
            .in2(_gnd_net_),
            .in3(N__5366),
            .lcout(\FSM_TEST_inst_slow.counter_idleZ0Z_1 ),
            .ltout(),
            .carryin(\FSM_TEST_inst_slow.counter_idle_cry_0 ),
            .carryout(\FSM_TEST_inst_slow.counter_idle_cry_1 ),
            .clk(N__10863),
            .ce(N__5549),
            .sr(N__10642));
    defparam \FSM_TEST_inst_slow.counter_idle_2_LC_10_18_2 .C_ON=1'b1;
    defparam \FSM_TEST_inst_slow.counter_idle_2_LC_10_18_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_idle_2_LC_10_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \FSM_TEST_inst_slow.counter_idle_2_LC_10_18_2  (
            .in0(N__5655),
            .in1(N__5525),
            .in2(_gnd_net_),
            .in3(N__5567),
            .lcout(\FSM_TEST_inst_slow.counter_idleZ0Z_2 ),
            .ltout(),
            .carryin(\FSM_TEST_inst_slow.counter_idle_cry_1 ),
            .carryout(\FSM_TEST_inst_slow.counter_idle_cry_2 ),
            .clk(N__10863),
            .ce(N__5549),
            .sr(N__10642));
    defparam \FSM_TEST_inst_slow.counter_idle_3_LC_10_18_3 .C_ON=1'b1;
    defparam \FSM_TEST_inst_slow.counter_idle_3_LC_10_18_3 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_idle_3_LC_10_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \FSM_TEST_inst_slow.counter_idle_3_LC_10_18_3  (
            .in0(N__5642),
            .in1(N__5606),
            .in2(_gnd_net_),
            .in3(N__5564),
            .lcout(\FSM_TEST_inst_slow.counter_idleZ0Z_3 ),
            .ltout(),
            .carryin(\FSM_TEST_inst_slow.counter_idle_cry_2 ),
            .carryout(\FSM_TEST_inst_slow.counter_idle_cry_3 ),
            .clk(N__10863),
            .ce(N__5549),
            .sr(N__10642));
    defparam \FSM_TEST_inst_slow.counter_idle_4_LC_10_18_4 .C_ON=1'b1;
    defparam \FSM_TEST_inst_slow.counter_idle_4_LC_10_18_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_idle_4_LC_10_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \FSM_TEST_inst_slow.counter_idle_4_LC_10_18_4  (
            .in0(N__5656),
            .in1(N__5624),
            .in2(_gnd_net_),
            .in3(N__5561),
            .lcout(\FSM_TEST_inst_slow.counter_idleZ0Z_4 ),
            .ltout(),
            .carryin(\FSM_TEST_inst_slow.counter_idle_cry_3 ),
            .carryout(\FSM_TEST_inst_slow.counter_idle_cry_4 ),
            .clk(N__10863),
            .ce(N__5549),
            .sr(N__10642));
    defparam \FSM_TEST_inst_slow.counter_idle_5_LC_10_18_5 .C_ON=1'b1;
    defparam \FSM_TEST_inst_slow.counter_idle_5_LC_10_18_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_idle_5_LC_10_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \FSM_TEST_inst_slow.counter_idle_5_LC_10_18_5  (
            .in0(N__5643),
            .in1(N__5509),
            .in2(_gnd_net_),
            .in3(N__5558),
            .lcout(\FSM_TEST_inst_slow.counter_idleZ0Z_5 ),
            .ltout(),
            .carryin(\FSM_TEST_inst_slow.counter_idle_cry_4 ),
            .carryout(\FSM_TEST_inst_slow.counter_idle_cry_5 ),
            .clk(N__10863),
            .ce(N__5549),
            .sr(N__10642));
    defparam \FSM_TEST_inst_slow.counter_idle_6_LC_10_18_6 .C_ON=1'b1;
    defparam \FSM_TEST_inst_slow.counter_idle_6_LC_10_18_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_idle_6_LC_10_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \FSM_TEST_inst_slow.counter_idle_6_LC_10_18_6  (
            .in0(N__5657),
            .in1(N__6180),
            .in2(_gnd_net_),
            .in3(N__5555),
            .lcout(\FSM_TEST_inst_slow.counter_idleZ0Z_6 ),
            .ltout(),
            .carryin(\FSM_TEST_inst_slow.counter_idle_cry_5 ),
            .carryout(\FSM_TEST_inst_slow.counter_idle_cry_6 ),
            .clk(N__10863),
            .ce(N__5549),
            .sr(N__10642));
    defparam \FSM_TEST_inst_slow.counter_idle_7_LC_10_18_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_idle_7_LC_10_18_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_idle_7_LC_10_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \FSM_TEST_inst_slow.counter_idle_7_LC_10_18_7  (
            .in0(N__5644),
            .in1(N__6212),
            .in2(_gnd_net_),
            .in3(N__5552),
            .lcout(\FSM_TEST_inst_slow.counter_idleZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10863),
            .ce(N__5549),
            .sr(N__10642));
    defparam \FSM_TEST_inst_slow.current_state_RNO_3_0_LC_10_19_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNO_3_0_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNO_3_0_LC_10_19_0 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNO_3_0_LC_10_19_0  (
            .in0(N__5536),
            .in1(N__5524),
            .in2(N__5513),
            .in3(N__5488),
            .lcout(\FSM_TEST_inst_slow.current_state_RNO_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.counter_din_RNO_0_3_LC_10_19_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_din_RNO_0_3_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.counter_din_RNO_0_3_LC_10_19_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \FSM_TEST_inst_slow.counter_din_RNO_0_3_LC_10_19_1  (
            .in0(N__5466),
            .in1(_gnd_net_),
            .in2(N__5450),
            .in3(N__6920),
            .lcout(\FSM_TEST_inst_slow.N_109_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.counter_din_RNID6M9_1_LC_10_19_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_din_RNID6M9_1_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.counter_din_RNID6M9_1_LC_10_19_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \FSM_TEST_inst_slow.counter_din_RNID6M9_1_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__5465),
            .in2(_gnd_net_),
            .in3(N__5445),
            .lcout(\FSM_TEST_inst_slow.N_106_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_4_0_LC_10_19_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_4_0_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_4_0_LC_10_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_RNO_4_0_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__5689),
            .in2(_gnd_net_),
            .in3(N__5749),
            .lcout(\FSM_TEST_inst_RAPIDA.G_24_0_a4_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.current_state_RNIV6JP_0_1_LC_10_19_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNIV6JP_0_1_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNIV6JP_0_1_LC_10_19_4 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNIV6JP_0_1_LC_10_19_4  (
            .in0(N__9003),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7850),
            .lcout(\FSM_TEST_inst_slow.current_state_d_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.current_state_RNIV6JP_1_LC_10_19_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNIV6JP_1_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNIV6JP_1_LC_10_19_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNIV6JP_1_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(N__7849),
            .in2(_gnd_net_),
            .in3(N__9002),
            .lcout(\FSM_TEST_inst_slow.N_134_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.current_state_RNO_5_0_LC_10_19_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNO_5_0_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNO_5_0_LC_10_19_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNO_5_0_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(N__5622),
            .in2(_gnd_net_),
            .in3(N__5604),
            .lcout(\FSM_TEST_inst_slow.current_state_RNO_5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_4_LC_10_20_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_4_LC_10_20_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_4_LC_10_20_0 .LUT_INIT=16'b0010011000101010;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_stat_4_LC_10_20_0  (
            .in0(N__6006),
            .in1(N__5720),
            .in2(N__6250),
            .in3(N__5588),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10876),
            .ce(),
            .sr(N__10634));
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_5_LC_10_20_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_5_LC_10_20_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_5_LC_10_20_1 .LUT_INIT=16'b0001111100100000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_stat_5_LC_10_20_1  (
            .in0(N__5582),
            .in1(N__6244),
            .in2(N__5726),
            .in3(N__5987),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10876),
            .ce(),
            .sr(N__10634));
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_3_LC_10_20_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_3_LC_10_20_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_3_LC_10_20_2 .LUT_INIT=16'b0000011010101010;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_stat_3_LC_10_20_2  (
            .in0(N__6984),
            .in1(N__5576),
            .in2(N__6249),
            .in3(N__5724),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10876),
            .ce(),
            .sr(N__10634));
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_RNIUUIP1_6_LC_10_20_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_RNIUUIP1_6_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_RNIUUIP1_6_LC_10_20_3 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_stat_RNIUUIP1_6_LC_10_20_3  (
            .in0(N__5984),
            .in1(N__6005),
            .in2(N__7017),
            .in3(N__6983),
            .lcout(),
            .ltout(\FSM_TEST_inst_RAPIDA.counter_statlde_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2_1_LC_10_20_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2_1_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2_1_LC_10_20_4 .LUT_INIT=16'b1100110001001100;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2_1_LC_10_20_4  (
            .in0(N__9412),
            .in1(N__11649),
            .in2(N__5570),
            .in3(N__11459),
            .lcout(\FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2Z0Z_1 ),
            .ltout(\FSM_TEST_inst_RAPIDA.current_state_fast_RNI571R2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_0_LC_10_20_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_0_LC_10_20_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_0_LC_10_20_5 .LUT_INIT=16'b0001111100100000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_stat_0_LC_10_20_5  (
            .in0(N__6616),
            .in1(N__6233),
            .in2(N__5753),
            .in3(N__5750),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10876),
            .ce(),
            .sr(N__10634));
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_1_LC_10_20_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_1_LC_10_20_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_1_LC_10_20_6 .LUT_INIT=16'b0011011100001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_stat_1_LC_10_20_6  (
            .in0(N__5732),
            .in1(N__5719),
            .in2(N__6248),
            .in3(N__5962),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10876),
            .ce(),
            .sr(N__10634));
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_2_LC_10_20_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_2_LC_10_20_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_stat_2_LC_10_20_7 .LUT_INIT=16'b0101011100100000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_stat_2_LC_10_20_7  (
            .in0(N__5718),
            .in1(N__6237),
            .in2(N__5699),
            .in3(N__5690),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_statZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10876),
            .ce(),
            .sr(N__10634));
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_c_0_LC_10_21_0 .C_ON=1'b1;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_c_0_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_c_0_LC_10_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_idle_cry_c_0_LC_10_21_0  (
            .in0(_gnd_net_),
            .in1(N__6417),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(\FSM_TEST_inst_RAPIDA.counter_idle_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_0_THRU_LUT4_0_LC_10_21_1 .C_ON=1'b1;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_0_THRU_LUT4_0_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_0_THRU_LUT4_0_LC_10_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_idle_cry_0_THRU_LUT4_0_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__6460),
            .in2(_gnd_net_),
            .in3(N__5672),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_idle_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\FSM_TEST_inst_RAPIDA.counter_idle_cry_0 ),
            .carryout(\FSM_TEST_inst_RAPIDA.counter_idle_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_1_THRU_LUT4_0_LC_10_21_2 .C_ON=1'b1;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_1_THRU_LUT4_0_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_1_THRU_LUT4_0_LC_10_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_idle_cry_1_THRU_LUT4_0_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__6439),
            .in2(_gnd_net_),
            .in3(N__5669),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_idle_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\FSM_TEST_inst_RAPIDA.counter_idle_cry_1 ),
            .carryout(\FSM_TEST_inst_RAPIDA.counter_idle_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_2_THRU_LUT4_0_LC_10_21_3 .C_ON=1'b1;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_2_THRU_LUT4_0_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_2_THRU_LUT4_0_LC_10_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_idle_cry_2_THRU_LUT4_0_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__6298),
            .in2(_gnd_net_),
            .in3(N__5666),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_idle_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\FSM_TEST_inst_RAPIDA.counter_idle_cry_2 ),
            .carryout(\FSM_TEST_inst_RAPIDA.counter_idle_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_3_THRU_LUT4_0_LC_10_21_4 .C_ON=1'b1;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_3_THRU_LUT4_0_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_cry_3_THRU_LUT4_0_LC_10_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_idle_cry_3_THRU_LUT4_0_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__6317),
            .in2(_gnd_net_),
            .in3(N__5663),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_idle_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\FSM_TEST_inst_RAPIDA.counter_idle_cry_3 ),
            .carryout(\FSM_TEST_inst_RAPIDA.counter_idle_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_5_LC_10_21_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_5_LC_10_21_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_5_LC_10_21_5 .LUT_INIT=16'b0001110001001100;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_idle_5_LC_10_21_5  (
            .in0(N__6484),
            .in1(N__6276),
            .in2(N__6528),
            .in3(N__5660),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10882),
            .ce(),
            .sr(N__10629));
    defparam \FSM_TEST_inst_RAPIDA.flag_input_reg_LC_10_22_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.flag_input_reg_LC_10_22_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.flag_input_reg_LC_10_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.flag_input_reg_LC_10_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6602),
            .lcout(\FSM_TEST_inst_RAPIDA.flag_input_regZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10888),
            .ce(),
            .sr(N__10624));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_13_LC_11_13_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_13_LC_11_13_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_13_LC_11_13_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_13_LC_11_13_7  (
            .in0(N__8980),
            .in1(N__6545),
            .in2(_gnd_net_),
            .in3(N__7827),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10823),
            .ce(N__7328),
            .sr(N__10662));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_1_LC_11_14_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_1_LC_11_14_0 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_1_LC_11_14_0 .LUT_INIT=16'b1111111110100101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_1_LC_11_14_0  (
            .in0(N__8956),
            .in1(_gnd_net_),
            .in2(N__7923),
            .in3(N__5786),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10827),
            .ce(N__7325),
            .sr(N__10657));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_82_LC_11_14_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_82_LC_11_14_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_82_LC_11_14_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_82_LC_11_14_1  (
            .in0(N__5780),
            .in1(N__7858),
            .in2(_gnd_net_),
            .in3(N__8958),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10827),
            .ce(N__7325),
            .sr(N__10657));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_0_LC_11_14_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_0_LC_11_14_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_0_LC_11_14_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_0_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__7851),
            .in2(_gnd_net_),
            .in3(N__8955),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10827),
            .ce(N__7325),
            .sr(N__10657));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_81_LC_11_14_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_81_LC_11_14_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_81_LC_11_14_4 .LUT_INIT=16'b1111111110100101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_81_LC_11_14_4  (
            .in0(N__8957),
            .in1(_gnd_net_),
            .in2(N__7924),
            .in3(N__5861),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10827),
            .ce(N__7325),
            .sr(N__10657));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_46_LC_11_15_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_46_LC_11_15_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_46_LC_11_15_1 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_46_LC_11_15_1  (
            .in0(N__8973),
            .in1(_gnd_net_),
            .in2(N__7901),
            .in3(N__5837),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10833),
            .ce(N__7321),
            .sr(N__10652));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_4_LC_11_15_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_4_LC_11_15_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_4_LC_11_15_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_4_LC_11_15_2  (
            .in0(N__5867),
            .in1(N__7766),
            .in2(_gnd_net_),
            .in3(N__8974),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10833),
            .ce(N__7321),
            .sr(N__10652));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_5_LC_11_15_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_5_LC_11_15_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_5_LC_11_15_3 .LUT_INIT=16'b1111111110100101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_5_LC_11_15_3  (
            .in0(N__8975),
            .in1(_gnd_net_),
            .in2(N__7902),
            .in3(N__5765),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10833),
            .ce(N__7321),
            .sr(N__10652));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_2_LC_11_15_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_2_LC_11_15_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_2_LC_11_15_4 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_2_LC_11_15_4  (
            .in0(N__5759),
            .in1(N__7761),
            .in2(_gnd_net_),
            .in3(N__8971),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10833),
            .ce(N__7321),
            .sr(N__10652));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_3_LC_11_15_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_3_LC_11_15_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_3_LC_11_15_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_3_LC_11_15_6  (
            .in0(N__5873),
            .in1(N__7762),
            .in2(_gnd_net_),
            .in3(N__8972),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10833),
            .ce(N__7321),
            .sr(N__10652));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_80_LC_11_15_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_80_LC_11_15_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_80_LC_11_15_7 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_80_LC_11_15_7  (
            .in0(N__8976),
            .in1(_gnd_net_),
            .in2(N__7903),
            .in3(N__5798),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10833),
            .ce(N__7321),
            .sr(N__10652));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_43_LC_11_16_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_43_LC_11_16_0 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_43_LC_11_16_0 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_43_LC_11_16_0  (
            .in0(N__5855),
            .in1(N__7561),
            .in2(_gnd_net_),
            .in3(N__8713),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10842),
            .ce(N__7318),
            .sr(N__10648));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_70_LC_11_16_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_70_LC_11_16_2 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_70_LC_11_16_2 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_70_LC_11_16_2  (
            .in0(N__6758),
            .in1(N__7563),
            .in2(_gnd_net_),
            .in3(N__8716),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10842),
            .ce(N__7318),
            .sr(N__10648));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_45_LC_11_16_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_45_LC_11_16_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_45_LC_11_16_3 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_45_LC_11_16_3  (
            .in0(N__8715),
            .in1(N__5810),
            .in2(_gnd_net_),
            .in3(N__7565),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10842),
            .ce(N__7318),
            .sr(N__10648));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_77_LC_11_16_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_77_LC_11_16_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_77_LC_11_16_4 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_77_LC_11_16_4  (
            .in0(N__5831),
            .in1(N__7564),
            .in2(_gnd_net_),
            .in3(N__8717),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10842),
            .ce(N__7318),
            .sr(N__10648));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_78_LC_11_16_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_78_LC_11_16_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_78_LC_11_16_5 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_78_LC_11_16_5  (
            .in0(N__8718),
            .in1(N__5822),
            .in2(_gnd_net_),
            .in3(N__7566),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10842),
            .ce(N__7318),
            .sr(N__10648));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_44_LC_11_16_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_44_LC_11_16_6 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_44_LC_11_16_6 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_44_LC_11_16_6  (
            .in0(N__5816),
            .in1(N__7562),
            .in2(_gnd_net_),
            .in3(N__8714),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10842),
            .ce(N__7318),
            .sr(N__10648));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_79_LC_11_16_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_79_LC_11_16_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_79_LC_11_16_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_79_LC_11_16_7  (
            .in0(N__8719),
            .in1(N__5804),
            .in2(_gnd_net_),
            .in3(N__7567),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10842),
            .ce(N__7318),
            .sr(N__10648));
    defparam \FSM_TEST_inst_slow.counter_stat_cry_c_0_LC_11_17_0 .C_ON=1'b1;
    defparam \FSM_TEST_inst_slow.counter_stat_cry_c_0_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.counter_stat_cry_c_0_LC_11_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \FSM_TEST_inst_slow.counter_stat_cry_c_0_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__6123),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\FSM_TEST_inst_slow.counter_stat_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.counter_stat_cry_0_THRU_LUT4_0_LC_11_17_1 .C_ON=1'b1;
    defparam \FSM_TEST_inst_slow.counter_stat_cry_0_THRU_LUT4_0_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.counter_stat_cry_0_THRU_LUT4_0_LC_11_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.counter_stat_cry_0_THRU_LUT4_0_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__6051),
            .in2(_gnd_net_),
            .in3(N__5930),
            .lcout(\FSM_TEST_inst_slow.counter_stat_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\FSM_TEST_inst_slow.counter_stat_cry_0 ),
            .carryout(\FSM_TEST_inst_slow.counter_stat_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.counter_stat_cry_1_THRU_LUT4_0_LC_11_17_2 .C_ON=1'b1;
    defparam \FSM_TEST_inst_slow.counter_stat_cry_1_THRU_LUT4_0_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.counter_stat_cry_1_THRU_LUT4_0_LC_11_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.counter_stat_cry_1_THRU_LUT4_0_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__6102),
            .in2(_gnd_net_),
            .in3(N__5927),
            .lcout(\FSM_TEST_inst_slow.counter_stat_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\FSM_TEST_inst_slow.counter_stat_cry_1 ),
            .carryout(\FSM_TEST_inst_slow.counter_stat_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.counter_stat_cry_2_THRU_LUT4_0_LC_11_17_3 .C_ON=1'b1;
    defparam \FSM_TEST_inst_slow.counter_stat_cry_2_THRU_LUT4_0_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.counter_stat_cry_2_THRU_LUT4_0_LC_11_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.counter_stat_cry_2_THRU_LUT4_0_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__6080),
            .in2(_gnd_net_),
            .in3(N__5924),
            .lcout(\FSM_TEST_inst_slow.counter_stat_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\FSM_TEST_inst_slow.counter_stat_cry_2 ),
            .carryout(\FSM_TEST_inst_slow.counter_stat_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.counter_stat_cry_3_THRU_LUT4_0_LC_11_17_4 .C_ON=1'b1;
    defparam \FSM_TEST_inst_slow.counter_stat_cry_3_THRU_LUT4_0_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.counter_stat_cry_3_THRU_LUT4_0_LC_11_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.counter_stat_cry_3_THRU_LUT4_0_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__6028),
            .in2(_gnd_net_),
            .in3(N__5921),
            .lcout(\FSM_TEST_inst_slow.counter_stat_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\FSM_TEST_inst_slow.counter_stat_cry_3 ),
            .carryout(\FSM_TEST_inst_slow.counter_stat_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.counter_stat_cry_4_THRU_LUT4_0_LC_11_17_5 .C_ON=1'b1;
    defparam \FSM_TEST_inst_slow.counter_stat_cry_4_THRU_LUT4_0_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.counter_stat_cry_4_THRU_LUT4_0_LC_11_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.counter_stat_cry_4_THRU_LUT4_0_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__9196),
            .in2(_gnd_net_),
            .in3(N__5918),
            .lcout(\FSM_TEST_inst_slow.counter_stat_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\FSM_TEST_inst_slow.counter_stat_cry_4 ),
            .carryout(\FSM_TEST_inst_slow.counter_stat_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.counter_stat_6_LC_11_17_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_stat_6_LC_11_17_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_stat_6_LC_11_17_6 .LUT_INIT=16'b0011010001110000;
    LogicCell40 \FSM_TEST_inst_slow.counter_stat_6_LC_11_17_6  (
            .in0(N__9250),
            .in1(N__9293),
            .in2(N__5911),
            .in3(N__5915),
            .lcout(\FSM_TEST_inst_slow.counter_statZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10850),
            .ce(),
            .sr(N__10643));
    defparam \FSM_TEST_inst_slow.current_state_RNO_6_0_LC_11_18_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNO_6_0_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNO_6_0_LC_11_18_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNO_6_0_LC_11_18_1  (
            .in0(N__6103),
            .in1(N__6078),
            .in2(N__5910),
            .in3(N__6124),
            .lcout(),
            .ltout(\FSM_TEST_inst_slow.current_state_ns_0_a3_1_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.current_state_RNO_1_0_LC_11_18_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNO_1_0_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNO_1_0_LC_11_18_2 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNO_1_0_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5882),
            .in3(N__5879),
            .lcout(\FSM_TEST_inst_slow.current_state_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.counter_stat_0_LC_11_18_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_stat_0_LC_11_18_3 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_stat_0_LC_11_18_3 .LUT_INIT=16'b0101011100100000;
    LogicCell40 \FSM_TEST_inst_slow.counter_stat_0_LC_11_18_3  (
            .in0(N__9287),
            .in1(N__9239),
            .in2(N__6617),
            .in3(N__6125),
            .lcout(\FSM_TEST_inst_slow.counter_statZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10857),
            .ce(),
            .sr(N__10638));
    defparam \FSM_TEST_inst_slow.counter_stat_2_LC_11_18_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_stat_2_LC_11_18_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_stat_2_LC_11_18_4 .LUT_INIT=16'b0000011011001100;
    LogicCell40 \FSM_TEST_inst_slow.counter_stat_2_LC_11_18_4  (
            .in0(N__6110),
            .in1(N__6104),
            .in2(N__9255),
            .in3(N__9291),
            .lcout(\FSM_TEST_inst_slow.counter_statZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10857),
            .ce(),
            .sr(N__10638));
    defparam \FSM_TEST_inst_slow.counter_stat_3_LC_11_18_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_stat_3_LC_11_18_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_stat_3_LC_11_18_5 .LUT_INIT=16'b0101011100100000;
    LogicCell40 \FSM_TEST_inst_slow.counter_stat_3_LC_11_18_5  (
            .in0(N__9288),
            .in1(N__9240),
            .in2(N__6089),
            .in3(N__6079),
            .lcout(\FSM_TEST_inst_slow.counter_statZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10857),
            .ce(),
            .sr(N__10638));
    defparam \FSM_TEST_inst_slow.counter_stat_1_LC_11_18_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_stat_1_LC_11_18_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_stat_1_LC_11_18_6 .LUT_INIT=16'b0011011100001000;
    LogicCell40 \FSM_TEST_inst_slow.counter_stat_1_LC_11_18_6  (
            .in0(N__6059),
            .in1(N__9290),
            .in2(N__9254),
            .in3(N__6053),
            .lcout(\FSM_TEST_inst_slow.counter_statZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10857),
            .ce(),
            .sr(N__10638));
    defparam \FSM_TEST_inst_slow.counter_stat_4_LC_11_18_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_stat_4_LC_11_18_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_stat_4_LC_11_18_7 .LUT_INIT=16'b0100011001001100;
    LogicCell40 \FSM_TEST_inst_slow.counter_stat_4_LC_11_18_7  (
            .in0(N__9289),
            .in1(N__6029),
            .in2(N__9259),
            .in3(N__6035),
            .lcout(\FSM_TEST_inst_slow.counter_statZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10857),
            .ce(),
            .sr(N__10638));
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_0_0_LC_11_19_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_0_0_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_0_0_LC_11_19_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_RNO_0_0_LC_11_19_0  (
            .in0(N__6008),
            .in1(N__5985),
            .in2(N__8463),
            .in3(N__5963),
            .lcout(\FSM_TEST_inst_RAPIDA.G_24_0_a4_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_RNI2J9G_LC_11_19_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_RNI2J9G_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_RNI2J9G_LC_11_19_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_RNI2J9G_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__8455),
            .in2(_gnd_net_),
            .in3(N__11193),
            .lcout(\FSM_TEST_inst_RAPIDA.N_126_1_i ),
            .ltout(\FSM_TEST_inst_RAPIDA.N_126_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_1_LC_11_19_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_1_LC_11_19_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_1_LC_11_19_2 .LUT_INIT=16'b0000011011001100;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_idle_1_LC_11_19_2  (
            .in0(N__5942),
            .in1(N__6459),
            .in2(N__5933),
            .in3(N__6520),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10864),
            .ce(),
            .sr(N__10635));
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_RNI2J9G_0_LC_11_19_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_RNI2J9G_0_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_RNI2J9G_0_LC_11_19_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_RNI2J9G_0_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__8454),
            .in2(_gnd_net_),
            .in3(N__11194),
            .lcout(\FSM_TEST_inst_RAPIDA.current_state_d_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.flag_output_1_LC_11_19_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.flag_output_1_LC_11_19_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.flag_output_1_LC_11_19_4 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.flag_output_1_LC_11_19_4  (
            .in0(N__11195),
            .in1(N__8462),
            .in2(N__11657),
            .in3(N__8061),
            .lcout(flag_signal),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10864),
            .ce(),
            .sr(N__10635));
    defparam \FSM_TEST_inst_slow.flag_input_reg_LC_11_19_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.flag_input_reg_LC_11_19_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.flag_input_reg_LC_11_19_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \FSM_TEST_inst_slow.flag_input_reg_LC_11_19_5  (
            .in0(N__8062),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\FSM_TEST_inst_slow.flag_input_regZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10864),
            .ce(),
            .sr(N__10635));
    defparam \FSM_TEST_inst_slow.current_state_RNO_4_0_LC_11_19_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNO_4_0_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNO_4_0_LC_11_19_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNO_4_0_LC_11_19_6  (
            .in0(N__7620),
            .in1(N__6210),
            .in2(N__6194),
            .in3(N__8768),
            .lcout(),
            .ltout(\FSM_TEST_inst_slow.current_state_RNO_4Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.current_state_RNO_0_0_LC_11_19_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNO_0_0_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNO_0_0_LC_11_19_7 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNO_0_0_LC_11_19_7  (
            .in0(N__6184),
            .in1(N__6158),
            .in2(N__6152),
            .in3(N__6149),
            .lcout(\FSM_TEST_inst_slow.N_134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_3_0_LC_11_20_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_3_0_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_3_0_LC_11_20_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_RNO_3_0_LC_11_20_0  (
            .in0(N__6335),
            .in1(N__11651),
            .in2(N__8468),
            .in3(N__6404),
            .lcout(\FSM_TEST_inst_RAPIDA.N_18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_0_LC_11_20_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_0_LC_11_20_1 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_0_LC_11_20_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_0_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__8467),
            .in2(_gnd_net_),
            .in3(N__11262),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10870),
            .ce(N__12152),
            .sr(N__10630));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_1_LC_11_20_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_1_LC_11_20_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_1_LC_11_20_2 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_1_LC_11_20_2  (
            .in0(N__11259),
            .in1(N__10330),
            .in2(_gnd_net_),
            .in3(N__6143),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10870),
            .ce(N__12152),
            .sr(N__10630));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_2_LC_11_20_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_2_LC_11_20_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_2_LC_11_20_3 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_2_LC_11_20_3  (
            .in0(N__11861),
            .in1(N__6137),
            .in2(_gnd_net_),
            .in3(N__11263),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10870),
            .ce(N__12152),
            .sr(N__10630));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_3_LC_11_20_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_3_LC_11_20_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_3_LC_11_20_4 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_3_LC_11_20_4  (
            .in0(N__11260),
            .in1(N__10331),
            .in2(_gnd_net_),
            .in3(N__6131),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10870),
            .ce(N__12152),
            .sr(N__10630));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_4_LC_11_20_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_4_LC_11_20_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_4_LC_11_20_5 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_4_LC_11_20_5  (
            .in0(N__10332),
            .in1(N__6365),
            .in2(_gnd_net_),
            .in3(N__11264),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10870),
            .ce(N__12152),
            .sr(N__10630));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_5_LC_11_20_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_5_LC_11_20_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_5_LC_11_20_6 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_5_LC_11_20_6  (
            .in0(N__11261),
            .in1(N__10333),
            .in2(_gnd_net_),
            .in3(N__6359),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10870),
            .ce(N__12152),
            .sr(N__10630));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_6_LC_11_20_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_6_LC_11_20_7 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_6_LC_11_20_7 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_6_LC_11_20_7  (
            .in0(N__11862),
            .in1(N__6353),
            .in2(_gnd_net_),
            .in3(N__11265),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10870),
            .ce(N__12152),
            .sr(N__10630));
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_4_LC_11_21_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_4_LC_11_21_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_4_LC_11_21_0 .LUT_INIT=16'b0001101000101010;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_idle_4_LC_11_21_0  (
            .in0(N__6316),
            .in1(N__6488),
            .in2(N__6530),
            .in3(N__6347),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10877),
            .ce(),
            .sr(N__10625));
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_6_0_LC_11_21_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_6_0_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_6_0_LC_11_21_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_RNO_6_0_LC_11_21_1  (
            .in0(N__6294),
            .in1(N__6315),
            .in2(N__6277),
            .in3(N__6341),
            .lcout(\FSM_TEST_inst_RAPIDA.G_24_0_a4_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_2_LC_11_21_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_2_LC_11_21_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_2_LC_11_21_2 .LUT_INIT=16'b0001111100100000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_idle_2_LC_11_21_2  (
            .in0(N__6329),
            .in1(N__6487),
            .in2(N__6529),
            .in3(N__6438),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10877),
            .ce(),
            .sr(N__10625));
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_3_LC_11_21_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_3_LC_11_21_3 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_3_LC_11_21_3 .LUT_INIT=16'b0011010001110000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_idle_3_LC_11_21_3  (
            .in0(N__6485),
            .in1(N__6521),
            .in2(N__6299),
            .in3(N__6323),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10877),
            .ce(),
            .sr(N__10625));
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_RNI23T81_5_LC_11_21_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_RNI23T81_5_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_RNI23T81_5_LC_11_21_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_idle_RNI23T81_5_LC_11_21_4  (
            .in0(N__6314),
            .in1(N__6293),
            .in2(N__6278),
            .in3(N__6434),
            .lcout(),
            .ltout(\FSM_TEST_inst_RAPIDA.counter_idlelde_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2_1_LC_11_21_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2_1_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2_1_LC_11_21_5 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2_1_LC_11_21_5  (
            .in0(N__11271),
            .in1(N__9420),
            .in2(N__6533),
            .in3(N__11650),
            .lcout(\FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1 ),
            .ltout(\FSM_TEST_inst_RAPIDA.current_state_fast_RNI9BBA2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_0_LC_11_21_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_0_LC_11_21_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_idle_0_LC_11_21_6 .LUT_INIT=16'b0000101001101010;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_idle_0_LC_11_21_6  (
            .in0(N__6419),
            .in1(N__6609),
            .in2(N__6491),
            .in3(N__6486),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_idleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10877),
            .ce(),
            .sr(N__10625));
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_7_0_LC_11_21_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_7_0_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_7_0_LC_11_21_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_RNO_7_0_LC_11_21_7  (
            .in0(N__11270),
            .in1(N__6461),
            .in2(N__6440),
            .in3(N__6418),
            .lcout(\FSM_TEST_inst_RAPIDA.G_24_0_a4_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_7_LC_11_22_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_7_LC_11_22_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_7_LC_11_22_0 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_7_LC_11_22_0  (
            .in0(N__11282),
            .in1(N__10340),
            .in2(_gnd_net_),
            .in3(N__6398),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10883),
            .ce(N__12151),
            .sr(N__10620));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_19_LC_11_22_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_19_LC_11_22_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_19_LC_11_22_1 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_19_LC_11_22_1  (
            .in0(N__10334),
            .in1(N__7112),
            .in2(_gnd_net_),
            .in3(N__11283),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10883),
            .ce(N__12151),
            .sr(N__10620));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_20_LC_11_22_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_20_LC_11_22_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_20_LC_11_22_2 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_20_LC_11_22_2  (
            .in0(N__11279),
            .in1(N__10335),
            .in2(_gnd_net_),
            .in3(N__6389),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10883),
            .ce(N__12151),
            .sr(N__10620));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_21_LC_11_22_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_21_LC_11_22_3 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_21_LC_11_22_3 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_21_LC_11_22_3  (
            .in0(N__10336),
            .in1(N__6383),
            .in2(_gnd_net_),
            .in3(N__11284),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10883),
            .ce(N__12151),
            .sr(N__10620));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_22_LC_11_22_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_22_LC_11_22_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_22_LC_11_22_4 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_22_LC_11_22_4  (
            .in0(N__11280),
            .in1(N__10337),
            .in2(_gnd_net_),
            .in3(N__6377),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10883),
            .ce(N__12151),
            .sr(N__10620));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_23_LC_11_22_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_23_LC_11_22_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_23_LC_11_22_6 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_23_LC_11_22_6  (
            .in0(N__11281),
            .in1(N__10338),
            .in2(_gnd_net_),
            .in3(N__6371),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10883),
            .ce(N__12151),
            .sr(N__10620));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_24_LC_11_22_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_24_LC_11_22_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_24_LC_11_22_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_24_LC_11_22_7  (
            .in0(N__10339),
            .in1(N__6623),
            .in2(_gnd_net_),
            .in3(N__11285),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10883),
            .ce(N__12151),
            .sr(N__10620));
    defparam CONSTANT_ONE_LUT4_LC_11_23_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_11_23_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_11_23_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_11_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_86_LC_12_11_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_86_LC_12_11_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_86_LC_12_11_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_86_LC_12_11_6  (
            .in0(N__6563),
            .in1(N__7811),
            .in2(_gnd_net_),
            .in3(N__9044),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10819),
            .ce(N__7334),
            .sr(N__10667));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_84_LC_12_12_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_84_LC_12_12_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_84_LC_12_12_4 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_84_LC_12_12_4  (
            .in0(N__6551),
            .in1(N__7807),
            .in2(_gnd_net_),
            .in3(N__9042),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10820),
            .ce(N__7333),
            .sr(N__10663));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_85_LC_12_12_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_85_LC_12_12_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_85_LC_12_12_5 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_85_LC_12_12_5  (
            .in0(N__9043),
            .in1(_gnd_net_),
            .in2(N__7915),
            .in3(N__6569),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10820),
            .ce(N__7333),
            .sr(N__10663));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_83_LC_12_13_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_83_LC_12_13_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_83_LC_12_13_0 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_83_LC_12_13_0  (
            .in0(N__8979),
            .in1(_gnd_net_),
            .in2(N__7914),
            .in3(N__6557),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10822),
            .ce(N__7332),
            .sr(N__10658));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_12_LC_12_13_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_12_LC_12_13_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_12_LC_12_13_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_12_LC_12_13_1  (
            .in0(N__6662),
            .in1(N__7800),
            .in2(_gnd_net_),
            .in3(N__8977),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10822),
            .ce(N__7332),
            .sr(N__10658));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_53_LC_12_13_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_53_LC_12_13_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_53_LC_12_13_6 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_53_LC_12_13_6  (
            .in0(N__8978),
            .in1(_gnd_net_),
            .in2(N__7913),
            .in3(N__6539),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10822),
            .ce(N__7332),
            .sr(N__10658));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_7_LC_12_14_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_7_LC_12_14_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_7_LC_12_14_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_7_LC_12_14_1  (
            .in0(N__6770),
            .in1(N__7781),
            .in2(_gnd_net_),
            .in3(N__8968),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10824),
            .ce(N__7329),
            .sr(N__10653));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_52_LC_12_14_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_52_LC_12_14_2 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_52_LC_12_14_2 .LUT_INIT=16'b1111111110100101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_52_LC_12_14_2  (
            .in0(N__8966),
            .in1(_gnd_net_),
            .in2(N__7904),
            .in3(N__6635),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10824),
            .ce(N__7329),
            .sr(N__10653));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_10_LC_12_14_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_10_LC_12_14_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_10_LC_12_14_3 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_10_LC_12_14_3  (
            .in0(N__6680),
            .in1(N__7773),
            .in2(_gnd_net_),
            .in3(N__8964),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10824),
            .ce(N__7329),
            .sr(N__10653));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_8_LC_12_14_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_8_LC_12_14_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_8_LC_12_14_4 .LUT_INIT=16'b1111111110100101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_8_LC_12_14_4  (
            .in0(N__8969),
            .in1(_gnd_net_),
            .in2(N__7906),
            .in3(N__6692),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10824),
            .ce(N__7329),
            .sr(N__10653));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_9_LC_12_14_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_9_LC_12_14_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_9_LC_12_14_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_9_LC_12_14_5  (
            .in0(N__6686),
            .in1(N__7785),
            .in2(_gnd_net_),
            .in3(N__8970),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10824),
            .ce(N__7329),
            .sr(N__10653));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_54_LC_12_14_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_54_LC_12_14_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_54_LC_12_14_6 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_54_LC_12_14_6  (
            .in0(N__8967),
            .in1(_gnd_net_),
            .in2(N__7905),
            .in3(N__6674),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10824),
            .ce(N__7329),
            .sr(N__10653));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_11_LC_12_14_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_11_LC_12_14_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_11_LC_12_14_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_11_LC_12_14_7  (
            .in0(N__6668),
            .in1(N__7774),
            .in2(_gnd_net_),
            .in3(N__8965),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10824),
            .ce(N__7329),
            .sr(N__10653));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_55_LC_12_15_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_55_LC_12_15_0 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_55_LC_12_15_0 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_55_LC_12_15_0  (
            .in0(N__6656),
            .in1(N__7753),
            .in2(_gnd_net_),
            .in3(N__8960),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10828),
            .ce(N__7326),
            .sr(N__10649));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_56_LC_12_15_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_56_LC_12_15_3 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_56_LC_12_15_3 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_56_LC_12_15_3  (
            .in0(N__8961),
            .in1(_gnd_net_),
            .in2(N__7899),
            .in3(N__6650),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10828),
            .ce(N__7326),
            .sr(N__10649));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_51_LC_12_15_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_51_LC_12_15_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_51_LC_12_15_4 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_51_LC_12_15_4  (
            .in0(N__6644),
            .in1(N__7752),
            .in2(_gnd_net_),
            .in3(N__8959),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10828),
            .ce(N__7326),
            .sr(N__10649));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_6_LC_12_15_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_6_LC_12_15_5 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_6_LC_12_15_5 .LUT_INIT=16'b1111111110100101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_6_LC_12_15_5  (
            .in0(N__8963),
            .in1(_gnd_net_),
            .in2(N__7900),
            .in3(N__6629),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10828),
            .ce(N__7326),
            .sr(N__10649));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_57_LC_12_15_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_57_LC_12_15_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_57_LC_12_15_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_57_LC_12_15_6  (
            .in0(N__6764),
            .in1(N__7757),
            .in2(_gnd_net_),
            .in3(N__8962),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10828),
            .ce(N__7326),
            .sr(N__10649));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_69_LC_12_16_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_69_LC_12_16_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_69_LC_12_16_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_69_LC_12_16_2  (
            .in0(N__6752),
            .in1(N__7536),
            .in2(_gnd_net_),
            .in3(N__8712),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10834),
            .ce(N__7322),
            .sr(N__10644));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_68_LC_12_16_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_68_LC_12_16_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_68_LC_12_16_4 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_68_LC_12_16_4  (
            .in0(N__6746),
            .in1(N__7535),
            .in2(_gnd_net_),
            .in3(N__8711),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10834),
            .ce(N__7322),
            .sr(N__10644));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_67_LC_12_16_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_67_LC_12_16_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_67_LC_12_16_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_67_LC_12_16_6  (
            .in0(N__7130),
            .in1(N__7534),
            .in2(_gnd_net_),
            .in3(N__8710),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10834),
            .ce(N__7322),
            .sr(N__10644));
    defparam \FSM_TEST_inst_slow.current_state_RNO_0_1_LC_12_17_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNO_0_1_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNO_0_1_LC_12_17_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNO_0_1_LC_12_17_0  (
            .in0(N__8651),
            .in1(N__6943),
            .in2(N__6916),
            .in3(N__6891),
            .lcout(\FSM_TEST_inst_slow.current_state_cnv_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.current_state_RNIV6JP_1_1_LC_12_17_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNIV6JP_1_1_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNIV6JP_1_1_LC_12_17_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNIV6JP_1_1_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__7457),
            .in2(_gnd_net_),
            .in3(N__8650),
            .lcout(\FSM_TEST_inst_slow.N_108_li ),
            .ltout(\FSM_TEST_inst_slow.N_108_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.current_state_RNIR2L81_0_1_LC_12_17_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNIR2L81_0_1_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNIR2L81_0_1_LC_12_17_2 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNIR2L81_0_1_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6740),
            .in3(N__7208),
            .lcout(\FSM_TEST_inst_slow.current_state_RNIR2L81_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.current_state_1_LC_12_17_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_1_LC_12_17_3 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.current_state_1_LC_12_17_3 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \FSM_TEST_inst_slow.current_state_1_LC_12_17_3  (
            .in0(N__7210),
            .in1(N__6725),
            .in2(_gnd_net_),
            .in3(N__7459),
            .lcout(\FSM_TEST_inst_slow.current_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10843),
            .ce(),
            .sr(N__10639));
    defparam \FSM_TEST_inst_slow.counter_din_2_LC_12_17_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_din_2_LC_12_17_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_din_2_LC_12_17_4 .LUT_INIT=16'b0110000010101010;
    LogicCell40 \FSM_TEST_inst_slow.counter_din_2_LC_12_17_4  (
            .in0(N__6912),
            .in1(N__6893),
            .in2(N__6716),
            .in3(N__7211),
            .lcout(\FSM_TEST_inst_slow.counter_dinZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10843),
            .ce(),
            .sr(N__10639));
    defparam \FSM_TEST_inst_slow.current_state_RNO_8_0_LC_12_17_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNO_8_0_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNO_8_0_LC_12_17_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNO_8_0_LC_12_17_5  (
            .in0(N__6944),
            .in1(N__6908),
            .in2(_gnd_net_),
            .in3(N__7458),
            .lcout(),
            .ltout(\FSM_TEST_inst_slow.current_state_RNO_8Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.current_state_RNO_2_0_LC_12_17_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_RNO_2_0_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.current_state_RNO_2_0_LC_12_17_6 .LUT_INIT=16'b0010101011111111;
    LogicCell40 \FSM_TEST_inst_slow.current_state_RNO_2_0_LC_12_17_6  (
            .in0(N__8652),
            .in1(N__6892),
            .in2(N__6875),
            .in3(N__7209),
            .lcout(),
            .ltout(\FSM_TEST_inst_slow.current_state_RNO_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.current_state_0_LC_12_17_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.current_state_0_LC_12_17_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.current_state_0_LC_12_17_7 .LUT_INIT=16'b1111110100001101;
    LogicCell40 \FSM_TEST_inst_slow.current_state_0_LC_12_17_7  (
            .in0(N__6872),
            .in1(N__6866),
            .in2(N__6857),
            .in3(N__8653),
            .lcout(\FSM_TEST_inst_slow.current_stateZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10843),
            .ce(),
            .sr(N__10639));
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNI9I121_8_LC_12_18_0 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNI9I121_8_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNI9I121_8_LC_12_18_0 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \config_register_latched_dec_inst.DYNCNF_1_RNI9I121_8_LC_12_18_0  (
            .in0(N__9536),
            .in1(N__6832),
            .in2(N__12083),
            .in3(N__10098),
            .lcout(s12_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \config_register_latched_dec_inst.DYNCNF_1_8_LC_12_18_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNCNF_1_8_LC_12_18_1 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNCNF_1_8_LC_12_18_1 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \config_register_latched_dec_inst.DYNCNF_1_8_LC_12_18_1  (
            .in0(N__9535),
            .in1(N__12063),
            .in2(N__6833),
            .in3(N__10085),
            .lcout(\config_register_latched_dec_inst.DYNCNF_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10851),
            .ce(N__8078),
            .sr(N__10636));
    defparam \config_register_latched_dec_inst.DYNCNF_1_9_LC_12_18_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNCNF_1_9_LC_12_18_2 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNCNF_1_9_LC_12_18_2 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \config_register_latched_dec_inst.DYNCNF_1_9_LC_12_18_2  (
            .in0(N__10086),
            .in1(N__9505),
            .in2(N__12082),
            .in3(N__6820),
            .lcout(\config_register_latched_dec_inst.DYNCNF_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10851),
            .ce(N__8078),
            .sr(N__10636));
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNIBK121_9_LC_12_18_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNIBK121_9_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNIBK121_9_LC_12_18_3 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \config_register_latched_dec_inst.DYNCNF_1_RNIBK121_9_LC_12_18_3  (
            .in0(N__6821),
            .in1(N__12070),
            .in2(N__9509),
            .in3(N__10088),
            .lcout(s13_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \config_register_latched_dec_inst.DYNCNF_1_0_LC_12_18_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNCNF_1_0_LC_12_18_4 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNCNF_1_0_LC_12_18_4 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \config_register_latched_dec_inst.DYNCNF_1_0_LC_12_18_4  (
            .in0(N__10087),
            .in1(N__8131),
            .in2(N__12081),
            .in3(N__6799),
            .lcout(\config_register_latched_dec_inst.DYNCNF_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10851),
            .ce(N__8078),
            .sr(N__10636));
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNIP1121_0_LC_12_18_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNIP1121_0_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNIP1121_0_LC_12_18_5 .LUT_INIT=16'b1010110010100000;
    LogicCell40 \config_register_latched_dec_inst.DYNCNF_1_RNIP1121_0_LC_12_18_5  (
            .in0(N__6800),
            .in1(N__12071),
            .in2(N__10105),
            .in3(N__8132),
            .lcout(\config_register_latched_dec_inst.DYNCNF_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \config_register_latched_dec_inst.DYNCNF_1_10_LC_12_18_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNCNF_1_10_LC_12_18_7 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNCNF_1_10_LC_12_18_7 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \config_register_latched_dec_inst.DYNCNF_1_10_LC_12_18_7  (
            .in0(N__8179),
            .in1(N__12062),
            .in2(N__8002),
            .in3(N__10084),
            .lcout(\config_register_latched_dec_inst.DYNCNF_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10851),
            .ce(N__8078),
            .sr(N__10636));
    defparam \FSM_TEST_inst_RAPIDA.counter_din_RNO_0_2_LC_12_19_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_din_RNO_0_2_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_din_RNO_0_2_LC_12_19_0 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_din_RNO_0_2_LC_12_19_0  (
            .in0(N__9932),
            .in1(N__9879),
            .in2(N__9977),
            .in3(N__11908),
            .lcout(),
            .ltout(\FSM_TEST_inst_RAPIDA.counter_din_3_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_din_2_LC_12_19_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_din_2_LC_12_19_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_din_2_LC_12_19_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_din_2_LC_12_19_1  (
            .in0(N__9971),
            .in1(N__8191),
            .in2(N__7040),
            .in3(N__11616),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_dinZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10858),
            .ce(),
            .sr(N__10631));
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_5_0_LC_12_19_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_5_0_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_5_0_LC_12_19_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_RNO_5_0_LC_12_19_2  (
            .in0(N__9931),
            .in1(N__9970),
            .in2(N__9909),
            .in3(N__9878),
            .lcout(),
            .ltout(\FSM_TEST_inst_RAPIDA.G_24_0_o4_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_2_0_LC_12_19_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_2_0_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_2_0_LC_12_19_3 .LUT_INIT=16'b1111101100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_RNO_2_0_LC_12_19_3  (
            .in0(N__8456),
            .in1(N__11613),
            .in2(N__7037),
            .in3(N__11220),
            .lcout(\FSM_TEST_inst_RAPIDA.N_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_1_0_LC_12_19_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_1_0_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_RNO_1_0_LC_12_19_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_RNO_1_0_LC_12_19_4  (
            .in0(N__11614),
            .in1(N__7034),
            .in2(N__7025),
            .in3(N__6992),
            .lcout(),
            .ltout(\FSM_TEST_inst_RAPIDA.G_24_0_a4_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.current_state_0_LC_12_19_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_0_LC_12_19_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.current_state_0_LC_12_19_5 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_0_LC_12_19_5  (
            .in0(N__6965),
            .in1(N__6959),
            .in2(N__6953),
            .in3(N__6950),
            .lcout(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10858),
            .ce(),
            .sr(N__10631));
    defparam \FSM_TEST_inst_RAPIDA.counter_din_1_LC_12_19_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_din_1_LC_12_19_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_din_1_LC_12_19_6 .LUT_INIT=16'b0111100001010000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_din_1_LC_12_19_6  (
            .in0(N__11615),
            .in1(N__9880),
            .in2(N__9940),
            .in3(N__11909),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_dinZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10858),
            .ce(),
            .sr(N__10631));
    defparam \FSM_TEST_inst_RAPIDA.counter_din_3_LC_12_19_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_din_3_LC_12_19_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_din_3_LC_12_19_7 .LUT_INIT=16'b0010100011110000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_din_3_LC_12_19_7  (
            .in0(N__11910),
            .in1(N__8192),
            .in2(N__9910),
            .in3(N__11617),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_dinZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10858),
            .ce(),
            .sr(N__10631));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_15_LC_12_20_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_15_LC_12_20_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_15_LC_12_20_0 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_15_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__11254),
            .in2(N__10341),
            .in3(N__7118),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10865),
            .ce(N__8233),
            .sr(N__10626));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_0_LC_12_20_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_0_LC_12_20_1 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_0_LC_12_20_1 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_0_LC_12_20_1  (
            .in0(N__11258),
            .in1(N__9413),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10865),
            .ce(N__8233),
            .sr(N__10626));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_5_LC_12_20_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_5_LC_12_20_2 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_5_LC_12_20_2 .LUT_INIT=16'b1111111111000011;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_5_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(N__11256),
            .in2(N__10342),
            .in3(N__7064),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10865),
            .ce(N__8233),
            .sr(N__10626));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_1_LC_12_20_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_1_LC_12_20_3 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_1_LC_12_20_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_1_LC_12_20_3  (
            .in0(N__7076),
            .in1(N__9414),
            .in2(_gnd_net_),
            .in3(N__11266),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10865),
            .ce(N__8233),
            .sr(N__10626));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_2_LC_12_20_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_2_LC_12_20_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_2_LC_12_20_4 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_2_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(N__11255),
            .in2(N__9424),
            .in3(N__7070),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10865),
            .ce(N__8233),
            .sr(N__10626));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_4_LC_12_20_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_4_LC_12_20_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_4_LC_12_20_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_4_LC_12_20_5  (
            .in0(N__7046),
            .in1(N__9419),
            .in2(_gnd_net_),
            .in3(N__11268),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10865),
            .ce(N__8233),
            .sr(N__10626));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_6_LC_12_20_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_6_LC_12_20_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_6_LC_12_20_6 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_6_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(N__11257),
            .in2(N__10343),
            .in3(N__7058),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10865),
            .ce(N__8233),
            .sr(N__10626));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_3_LC_12_20_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_3_LC_12_20_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_3_LC_12_20_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_3_LC_12_20_7  (
            .in0(N__7052),
            .in1(N__9418),
            .in2(_gnd_net_),
            .in3(N__11267),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10865),
            .ce(N__8233),
            .sr(N__10626));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_13_LC_12_21_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_13_LC_12_21_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_13_LC_12_21_4 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_13_LC_12_21_4  (
            .in0(N__10324),
            .in1(N__8243),
            .in2(_gnd_net_),
            .in3(N__11286),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10871),
            .ce(N__8237),
            .sr(N__10621));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_14_LC_12_21_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_14_LC_12_21_6 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_14_LC_12_21_6 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_14_LC_12_21_6  (
            .in0(N__10325),
            .in1(N__7124),
            .in2(_gnd_net_),
            .in3(N__11287),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10871),
            .ce(N__8237),
            .sr(N__10621));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_18_LC_12_22_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_18_LC_12_22_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_18_LC_12_22_0 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_18_LC_12_22_0  (
            .in0(N__10326),
            .in1(N__9755),
            .in2(_gnd_net_),
            .in3(N__11275),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10878),
            .ce(N__12149),
            .sr(N__10615));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_79_LC_12_22_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_79_LC_12_22_2 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_79_LC_12_22_2 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_79_LC_12_22_2  (
            .in0(N__11045),
            .in1(N__7100),
            .in2(_gnd_net_),
            .in3(N__11278),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10878),
            .ce(N__12149),
            .sr(N__10615));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_27_LC_12_22_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_27_LC_12_22_3 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_27_LC_12_22_3 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_27_LC_12_22_3  (
            .in0(N__11273),
            .in1(N__10328),
            .in2(_gnd_net_),
            .in3(N__7082),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10878),
            .ce(N__12149),
            .sr(N__10615));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_25_LC_12_22_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_25_LC_12_22_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_25_LC_12_22_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_25_LC_12_22_4  (
            .in0(N__7106),
            .in1(N__10329),
            .in2(_gnd_net_),
            .in3(N__11276),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10878),
            .ce(N__12149),
            .sr(N__10615));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_78_LC_12_22_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_78_LC_12_22_5 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_78_LC_12_22_5 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_78_LC_12_22_5  (
            .in0(N__11274),
            .in1(N__11044),
            .in2(_gnd_net_),
            .in3(N__7094),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10878),
            .ce(N__12149),
            .sr(N__10615));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_77_LC_12_22_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_77_LC_12_22_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_77_LC_12_22_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_77_LC_12_22_6  (
            .in0(N__11864),
            .in1(N__8408),
            .in2(_gnd_net_),
            .in3(N__11277),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10878),
            .ce(N__12149),
            .sr(N__10615));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_26_LC_12_22_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_26_LC_12_22_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_26_LC_12_22_7 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_26_LC_12_22_7  (
            .in0(N__11272),
            .in1(N__10327),
            .in2(_gnd_net_),
            .in3(N__7088),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10878),
            .ce(N__12149),
            .sr(N__10615));
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_4_0_LC_12_23_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_4_0_LC_12_23_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_4_0_LC_12_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.CLK_uC_4_0_LC_12_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7184),
            .lcout(\FSM_TEST_inst_RAPIDA.CLK_uC_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10884),
            .ce(),
            .sr(N__10611));
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_6_0_LC_12_23_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_6_0_LC_12_23_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_6_0_LC_12_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.CLK_uC_6_0_LC_12_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7172),
            .lcout(\FSM_TEST_inst_RAPIDA.CLK_uC_6Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10884),
            .ce(),
            .sr(N__10611));
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_3_0_LC_12_23_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_3_0_LC_12_23_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_3_0_LC_12_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.CLK_uC_3_0_LC_12_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8396),
            .lcout(\FSM_TEST_inst_RAPIDA.CLK_uC_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10884),
            .ce(),
            .sr(N__10611));
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_5_0_LC_12_23_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_5_0_LC_12_23_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_5_0_LC_12_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.CLK_uC_5_0_LC_12_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7178),
            .lcout(\FSM_TEST_inst_RAPIDA.CLK_uC_5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10884),
            .ce(),
            .sr(N__10611));
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_6b_0_LC_12_23_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_6b_0_LC_12_23_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_6b_0_LC_12_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.CLK_uC_6b_0_LC_12_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7166),
            .lcout(\FSM_TEST_inst_RAPIDA.CLK_uC_6bZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10884),
            .ce(),
            .sr(N__10611));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_61_LC_13_15_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_61_LC_13_15_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_61_LC_13_15_3 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_61_LC_13_15_3  (
            .in0(N__8941),
            .in1(N__7154),
            .in2(_gnd_net_),
            .in3(N__7799),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10825),
            .ce(N__7330),
            .sr(N__10645));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_58_LC_13_15_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_58_LC_13_15_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_58_LC_13_15_4 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_58_LC_13_15_4  (
            .in0(N__7796),
            .in1(N__7160),
            .in2(_gnd_net_),
            .in3(N__8938),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10825),
            .ce(N__7330),
            .sr(N__10645));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_60_LC_13_15_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_60_LC_13_15_5 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_60_LC_13_15_5 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_60_LC_13_15_5  (
            .in0(N__8940),
            .in1(N__7142),
            .in2(_gnd_net_),
            .in3(N__7798),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10825),
            .ce(N__7330),
            .sr(N__10645));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_59_LC_13_15_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_59_LC_13_15_7 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_59_LC_13_15_7 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_59_LC_13_15_7  (
            .in0(N__8939),
            .in1(N__7148),
            .in2(_gnd_net_),
            .in3(N__7797),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10825),
            .ce(N__7330),
            .sr(N__10645));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_62_LC_13_16_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_62_LC_13_16_0 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_62_LC_13_16_0 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_62_LC_13_16_0  (
            .in0(N__7136),
            .in1(N__7568),
            .in2(_gnd_net_),
            .in3(N__8720),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10829),
            .ce(N__7327),
            .sr(N__10640));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_66_LC_13_16_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_66_LC_13_16_1 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_66_LC_13_16_1 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_66_LC_13_16_1  (
            .in0(N__8724),
            .in1(N__7952),
            .in2(_gnd_net_),
            .in3(N__7572),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10829),
            .ce(N__7327),
            .sr(N__10640));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_64_LC_13_16_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_64_LC_13_16_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_64_LC_13_16_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_64_LC_13_16_2  (
            .in0(N__7340),
            .in1(N__7569),
            .in2(_gnd_net_),
            .in3(N__8722),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10829),
            .ce(N__7327),
            .sr(N__10640));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_65_LC_13_16_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_65_LC_13_16_5 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_65_LC_13_16_5 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_65_LC_13_16_5  (
            .in0(N__8723),
            .in1(N__7958),
            .in2(_gnd_net_),
            .in3(N__7571),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10829),
            .ce(N__7327),
            .sr(N__10640));
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_63_LC_13_16_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_63_LC_13_16_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.bit_sequence_stat_63_LC_13_16_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_slow.bit_sequence_stat_63_LC_13_16_7  (
            .in0(N__8721),
            .in1(N__7946),
            .in2(_gnd_net_),
            .in3(N__7570),
            .lcout(\FSM_TEST_inst_slow.bit_sequence_statZ0Z_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10829),
            .ce(N__7327),
            .sr(N__10640));
    defparam \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5D1_0_LC_13_17_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5D1_0_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5D1_0_LC_13_17_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5D1_0_LC_13_17_0  (
            .in0(N__11598),
            .in1(N__8496),
            .in2(N__9085),
            .in3(N__11269),
            .lcout(N_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divisor_inst_2.counter_RNIFD27_2_LC_13_17_1 .C_ON=1'b0;
    defparam \divisor_inst_2.counter_RNIFD27_2_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \divisor_inst_2.counter_RNIFD27_2_LC_13_17_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \divisor_inst_2.counter_RNIFD27_2_LC_13_17_1  (
            .in0(N__9163),
            .in1(_gnd_net_),
            .in2(N__9110),
            .in3(N__9130),
            .lcout(counter_RNIFD27_2),
            .ltout(counter_RNIFD27_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_slow.SEL_0_RNI25J31_LC_13_17_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.SEL_0_RNI25J31_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_slow.SEL_0_RNI25J31_LC_13_17_2 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \FSM_TEST_inst_slow.SEL_0_RNI25J31_LC_13_17_2  (
            .in0(N__8534),
            .in1(N__8513),
            .in2(N__7253),
            .in3(N__8709),
            .lcout(N_3_0),
            .ltout(N_3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \config_register_latched_dec_inst.STATCNF_1_RNO_0_LC_13_17_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.STATCNF_1_RNO_0_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst.STATCNF_1_RNO_0_LC_13_17_3 .LUT_INIT=16'b0000110000111111;
    LogicCell40 \config_register_latched_dec_inst.STATCNF_1_RNO_0_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__8351),
            .in2(N__7250),
            .in3(N__7247),
            .lcout(\config_register_latched_dec_inst.N_378_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divisor_inst_2.counter_RNISR1F_2_LC_13_17_5 .C_ON=1'b0;
    defparam \divisor_inst_2.counter_RNISR1F_2_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \divisor_inst_2.counter_RNISR1F_2_LC_13_17_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \divisor_inst_2.counter_RNISR1F_2_LC_13_17_5  (
            .in0(N__9162),
            .in1(N__9129),
            .in2(N__9109),
            .in3(N__8533),
            .lcout(counter_RNISR1F_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divisor_inst_2.clk_out_LC_13_17_6 .C_ON=1'b0;
    defparam \divisor_inst_2.clk_out_LC_13_17_6 .SEQ_MODE=4'b1010;
    defparam \divisor_inst_2.clk_out_LC_13_17_6 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \divisor_inst_2.clk_out_LC_13_17_6  (
            .in0(N__8535),
            .in1(N__9164),
            .in2(N__9139),
            .in3(N__9107),
            .lcout(clk_continuous_slow),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10835),
            .ce(),
            .sr(N__10637));
    defparam \FSM_TEST_inst_RAPIDA.MOSI_er_LC_13_18_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.MOSI_er_LC_13_18_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.MOSI_er_LC_13_18_0 .LUT_INIT=16'b0101000010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.MOSI_er_LC_13_18_0  (
            .in0(N__11149),
            .in1(N__8099),
            .in2(N__9671),
            .in3(N__8433),
            .lcout(mosi_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10844),
            .ce(N__11642),
            .sr(N__10632));
    defparam \divisor_inst.clk_out_RNI3LEM_LC_13_18_1 .C_ON=1'b0;
    defparam \divisor_inst.clk_out_RNI3LEM_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \divisor_inst.clk_out_RNI3LEM_LC_13_18_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \divisor_inst.clk_out_RNI3LEM_LC_13_18_1  (
            .in0(N__11992),
            .in1(N__11930),
            .in2(_gnd_net_),
            .in3(N__11960),
            .lcout(clk_out_RNI3LEM),
            .ltout(clk_out_RNI3LEM_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.flag_output_1_RNIVLAE1_LC_13_18_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.flag_output_1_RNIVLAE1_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.flag_output_1_RNIVLAE1_LC_13_18_2 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \FSM_TEST_inst_RAPIDA.flag_output_1_RNIVLAE1_LC_13_18_2  (
            .in0(N__11148),
            .in1(N__8068),
            .in2(N__8087),
            .in3(N__8432),
            .lcout(N_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIHTFF_1_LC_13_18_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIHTFF_1_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIHTFF_1_LC_13_18_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIHTFF_1_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(N__8486),
            .in2(_gnd_net_),
            .in3(N__11147),
            .lcout(\FSM_TEST_inst_RAPIDA.N_100_li ),
            .ltout(\FSM_TEST_inst_RAPIDA.N_100_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5D1_LC_13_18_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5D1_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5D1_LC_13_18_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5D1_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(N__9081),
            .in2(N__8084),
            .in3(N__11599),
            .lcout(\FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5DZ0Z1 ),
            .ltout(\FSM_TEST_inst_RAPIDA.SEL_0_RNI7M5DZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.SEL_0_RNI8H3V3_LC_13_18_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.SEL_0_RNI8H3V3_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.SEL_0_RNI8H3V3_LC_13_18_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.SEL_0_RNI8H3V3_LC_13_18_5  (
            .in0(N__8365),
            .in1(_gnd_net_),
            .in2(N__8081),
            .in3(N__8350),
            .lcout(N_378_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mosi_output_obuf_RNO_LC_13_18_7.C_ON=1'b0;
    defparam mosi_output_obuf_RNO_LC_13_18_7.SEQ_MODE=4'b0000;
    defparam mosi_output_obuf_RNO_LC_13_18_7.LUT_INIT=16'b1110111001000100;
    LogicCell40 mosi_output_obuf_RNO_LC_13_18_7 (
            .in0(N__8069),
            .in1(N__8045),
            .in2(_gnd_net_),
            .in3(N__8039),
            .lcout(mosi_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNIR83V_10_LC_13_19_0 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNIR83V_10_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst.DYNCNF_1_RNIR83V_10_LC_13_19_0 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \config_register_latched_dec_inst.DYNCNF_1_RNIR83V_10_LC_13_19_0  (
            .in0(N__10082),
            .in1(N__12095),
            .in2(N__8180),
            .in3(N__8003),
            .lcout(s14_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \config_register_latched_dec_inst.STATCNF_1_0_LC_13_19_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.STATCNF_1_0_LC_13_19_2 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.STATCNF_1_0_LC_13_19_2 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \config_register_latched_dec_inst.STATCNF_1_0_LC_13_19_2  (
            .in0(N__10081),
            .in1(N__12096),
            .in2(N__10153),
            .in3(N__10123),
            .lcout(\config_register_latched_dec_inst.STATCNF_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10852),
            .ce(N__7967),
            .sr(N__10627));
    defparam flag_output_0_ret_RNI1E8N2_LC_13_19_5.C_ON=1'b0;
    defparam flag_output_0_ret_RNI1E8N2_LC_13_19_5.SEQ_MODE=4'b0000;
    defparam flag_output_0_ret_RNI1E8N2_LC_13_19_5.LUT_INIT=16'b0010001000110000;
    LogicCell40 flag_output_0_ret_RNI1E8N2_LC_13_19_5 (
            .in0(N__9343),
            .in1(N__8290),
            .in2(N__8326),
            .in3(N__8352),
            .lcout(flag_output_0_ret_RNI1E8NZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_din_RNI9NO1_1_LC_13_19_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_din_RNI9NO1_1_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_din_RNI9NO1_1_LC_13_19_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_din_RNI9NO1_1_LC_13_19_6  (
            .in0(N__9973),
            .in1(N__9936),
            .in2(_gnd_net_),
            .in3(N__9873),
            .lcout(\FSM_TEST_inst_RAPIDA.N_101_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_RNI78E11_1_LC_13_19_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_RNI78E11_1_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_RNI78E11_1_LC_13_19_7 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_fast_RNI78E11_1_LC_13_19_7  (
            .in0(N__9387),
            .in1(N__11618),
            .in2(_gnd_net_),
            .in3(N__11219),
            .lcout(\FSM_TEST_inst_RAPIDA.current_state_fast_RNI78E11Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \config_register_latched_dec_inst.DYNSR_10_LC_13_20_0 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNSR_10_LC_13_20_0 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNSR_10_LC_13_20_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \config_register_latched_dec_inst.DYNSR_10_LC_13_20_0  (
            .in0(N__10083),
            .in1(N__8175),
            .in2(_gnd_net_),
            .in3(N__9499),
            .lcout(\config_register_latched_dec_inst.DYNSRZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10859),
            .ce(N__9478),
            .sr(N__10622));
    defparam \config_register_latched_dec_inst.STATSR_0_LC_13_20_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.STATSR_0_LC_13_20_3 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.STATSR_0_LC_13_20_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \config_register_latched_dec_inst.STATSR_0_LC_13_20_3  (
            .in0(N__10079),
            .in1(N__8156),
            .in2(_gnd_net_),
            .in3(N__10149),
            .lcout(\config_register_latched_dec_inst.STATSRZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10859),
            .ce(N__9478),
            .sr(N__10622));
    defparam \config_register_latched_dec_inst.DYNSR_1_LC_13_20_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNSR_1_LC_13_20_6 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNSR_1_LC_13_20_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \config_register_latched_dec_inst.DYNSR_1_LC_13_20_6  (
            .in0(N__8123),
            .in1(N__10080),
            .in2(_gnd_net_),
            .in3(N__9314),
            .lcout(\config_register_latched_dec_inst.DYNSRZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10859),
            .ce(N__9478),
            .sr(N__10622));
    defparam \config_register_latched_dec_inst.DYNSR_0_LC_13_20_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNSR_0_LC_13_20_7 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNSR_0_LC_13_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \config_register_latched_dec_inst.DYNSR_0_LC_13_20_7  (
            .in0(N__10078),
            .in1(N__8155),
            .in2(_gnd_net_),
            .in3(N__8124),
            .lcout(\config_register_latched_dec_inst.DYNSRZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10859),
            .ce(N__9478),
            .sr(N__10622));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_10_LC_13_21_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_10_LC_13_21_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_10_LC_13_21_0 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_10_LC_13_21_0  (
            .in0(N__11481),
            .in1(N__8255),
            .in2(_gnd_net_),
            .in3(N__10245),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10866),
            .ce(N__8232),
            .sr(N__10616));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_11_LC_13_21_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_11_LC_13_21_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_11_LC_13_21_1 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_11_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(N__11477),
            .in2(N__10311),
            .in3(N__8105),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10866),
            .ce(N__8232),
            .sr(N__10616));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_8_LC_13_21_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_8_LC_13_21_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_8_LC_13_21_3 .LUT_INIT=16'b1111111111000011;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_8_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(N__11480),
            .in2(N__10314),
            .in3(N__8267),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10866),
            .ce(N__8232),
            .sr(N__10616));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_7_LC_13_21_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_7_LC_13_21_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_7_LC_13_21_5 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_7_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(N__11479),
            .in2(N__10313),
            .in3(N__8273),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10866),
            .ce(N__8232),
            .sr(N__10616));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_9_LC_13_21_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_9_LC_13_21_6 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_9_LC_13_21_6 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_9_LC_13_21_6  (
            .in0(N__11482),
            .in1(N__8261),
            .in2(_gnd_net_),
            .in3(N__10258),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10866),
            .ce(N__8232),
            .sr(N__10616));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_12_LC_13_21_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_12_LC_13_21_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_din_12_LC_13_21_7 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_din_12_LC_13_21_7  (
            .in0(_gnd_net_),
            .in1(N__11478),
            .in2(N__10312),
            .in3(N__8249),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_dinZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10866),
            .ce(N__8232),
            .sr(N__10616));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_59_LC_13_22_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_59_LC_13_22_0 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_59_LC_13_22_0 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_59_LC_13_22_0  (
            .in0(N__11041),
            .in1(N__9608),
            .in2(_gnd_net_),
            .in3(N__11488),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10872),
            .ce(N__12146),
            .sr(N__10612));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_54_LC_13_22_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_54_LC_13_22_1 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_54_LC_13_22_1 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_54_LC_13_22_1  (
            .in0(N__11483),
            .in1(N__11040),
            .in2(_gnd_net_),
            .in3(N__9443),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10872),
            .ce(N__12146),
            .sr(N__10612));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_29_LC_13_22_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_29_LC_13_22_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_29_LC_13_22_2 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_29_LC_13_22_2  (
            .in0(N__10259),
            .in1(N__8204),
            .in2(_gnd_net_),
            .in3(N__11487),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10872),
            .ce(N__12146),
            .sr(N__10612));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_28_LC_13_22_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_28_LC_13_22_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_28_LC_13_22_4 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_28_LC_13_22_4  (
            .in0(N__11039),
            .in1(N__8210),
            .in2(_gnd_net_),
            .in3(N__11486),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10872),
            .ce(N__12146),
            .sr(N__10612));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_60_LC_13_22_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_60_LC_13_22_5 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_60_LC_13_22_5 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_60_LC_13_22_5  (
            .in0(N__11485),
            .in1(N__11042),
            .in2(_gnd_net_),
            .in3(N__8198),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10872),
            .ce(N__12146),
            .sr(N__10612));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_76_LC_13_22_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_76_LC_13_22_6 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_76_LC_13_22_6 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_76_LC_13_22_6  (
            .in0(N__11043),
            .in1(N__9620),
            .in2(_gnd_net_),
            .in3(N__11489),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10872),
            .ce(N__12146),
            .sr(N__10612));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_55_LC_13_22_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_55_LC_13_22_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_55_LC_13_22_7 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_55_LC_13_22_7  (
            .in0(N__11484),
            .in1(N__11863),
            .in2(_gnd_net_),
            .in3(N__8402),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10872),
            .ce(N__12146),
            .sr(N__10612));
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_2_0_LC_13_23_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_2_0_LC_13_23_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_2_0_LC_13_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.CLK_uC_2_0_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8383),
            .lcout(\FSM_TEST_inst_RAPIDA.CLK_uC_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10879),
            .ce(),
            .sr(N__10608));
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_6c_0_LC_13_23_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_6c_0_LC_13_23_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_6c_0_LC_13_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.CLK_uC_6c_0_LC_13_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8390),
            .lcout(CLK_uC_6c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10879),
            .ce(),
            .sr(N__10608));
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_LC_13_23_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_LC_13_23_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.CLK_uC_LC_13_23_7 .LUT_INIT=16'b1111011010010000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.CLK_uC_LC_13_23_7  (
            .in0(N__11466),
            .in1(N__9425),
            .in2(N__8384),
            .in3(N__11972),
            .lcout(\FSM_TEST_inst_RAPIDA.CLK_uCZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10879),
            .ce(),
            .sr(N__10608));
    defparam flag_output_ret_LC_14_17_1.C_ON=1'b0;
    defparam flag_output_ret_LC_14_17_1.SEQ_MODE=4'b1010;
    defparam flag_output_ret_LC_14_17_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 flag_output_ret_LC_14_17_1 (
            .in0(N__8372),
            .in1(N__8366),
            .in2(_gnd_net_),
            .in3(N__8353),
            .lcout(sel_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10830),
            .ce(),
            .sr(N__10633));
    defparam flag_output_0_ret_LC_14_17_2.C_ON=1'b0;
    defparam flag_output_0_ret_LC_14_17_2.SEQ_MODE=4'b1010;
    defparam flag_output_0_ret_LC_14_17_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 flag_output_0_ret_LC_14_17_2 (
            .in0(N__8354),
            .in1(N__9347),
            .in2(_gnd_net_),
            .in3(N__8327),
            .lcout(clk_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10830),
            .ce(),
            .sr(N__10633));
    defparam \divisor_inst_2.counter_1_LC_14_17_3 .C_ON=1'b0;
    defparam \divisor_inst_2.counter_1_LC_14_17_3 .SEQ_MODE=4'b1010;
    defparam \divisor_inst_2.counter_1_LC_14_17_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \divisor_inst_2.counter_1_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__9134),
            .in2(_gnd_net_),
            .in3(N__9160),
            .lcout(\divisor_inst_2.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10830),
            .ce(),
            .sr(N__10633));
    defparam \divisor_inst_2.counter_0_LC_14_17_4 .C_ON=1'b0;
    defparam \divisor_inst_2.counter_0_LC_14_17_4 .SEQ_MODE=4'b1010;
    defparam \divisor_inst_2.counter_0_LC_14_17_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \divisor_inst_2.counter_0_LC_14_17_4  (
            .in0(N__9135),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\divisor_inst_2.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10830),
            .ce(),
            .sr(N__10633));
    defparam \FSM_TEST_inst_slow.counter_stat_5_LC_14_17_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.counter_stat_5_LC_14_17_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.counter_stat_5_LC_14_17_5 .LUT_INIT=16'b0100011001001100;
    LogicCell40 \FSM_TEST_inst_slow.counter_stat_5_LC_14_17_5  (
            .in0(N__9292),
            .in1(N__9182),
            .in2(N__9260),
            .in3(N__9206),
            .lcout(\FSM_TEST_inst_slow.counter_statZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10830),
            .ce(),
            .sr(N__10633));
    defparam \divisor_inst_2.counter_2_LC_14_17_6 .C_ON=1'b0;
    defparam \divisor_inst_2.counter_2_LC_14_17_6 .SEQ_MODE=4'b1010;
    defparam \divisor_inst_2.counter_2_LC_14_17_6 .LUT_INIT=16'b0110110001101100;
    LogicCell40 \divisor_inst_2.counter_2_LC_14_17_6  (
            .in0(N__9161),
            .in1(N__9108),
            .in2(N__9140),
            .in3(_gnd_net_),
            .lcout(\divisor_inst_2.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10830),
            .ce(),
            .sr(N__10633));
    defparam \FSM_TEST_inst_RAPIDA.SEL_0_LC_14_17_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.SEL_0_LC_14_17_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.SEL_0_LC_14_17_7 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.SEL_0_LC_14_17_7  (
            .in0(N__8497),
            .in1(N__11619),
            .in2(N__9086),
            .in3(N__11534),
            .lcout(\FSM_TEST_inst_RAPIDA.aux_selection_fast_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10830),
            .ce(),
            .sr(N__10633));
    defparam \FSM_TEST_inst_slow.SEL_0_LC_14_18_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.SEL_0_LC_14_18_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.SEL_0_LC_14_18_2 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \FSM_TEST_inst_slow.SEL_0_LC_14_18_2  (
            .in0(N__8512),
            .in1(N__9012),
            .in2(N__8555),
            .in3(N__8536),
            .lcout(\FSM_TEST_inst_slow.aux_selection_slow_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10836),
            .ce(),
            .sr(N__10628));
    defparam \divisor_inst.clk_out_LC_14_18_3 .C_ON=1'b0;
    defparam \divisor_inst.clk_out_LC_14_18_3 .SEQ_MODE=4'b1010;
    defparam \divisor_inst.clk_out_LC_14_18_3 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \divisor_inst.clk_out_LC_14_18_3  (
            .in0(N__11935),
            .in1(N__11998),
            .in2(_gnd_net_),
            .in3(N__11964),
            .lcout(clk_continuous_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10836),
            .ce(),
            .sr(N__10628));
    defparam \divisor_inst.counter_1_LC_14_18_4 .C_ON=1'b0;
    defparam \divisor_inst.counter_1_LC_14_18_4 .SEQ_MODE=4'b1010;
    defparam \divisor_inst.counter_1_LC_14_18_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \divisor_inst.counter_1_LC_14_18_4  (
            .in0(N__11997),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11934),
            .lcout(divisor_inst_counter_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10836),
            .ce(),
            .sr(N__10628));
    defparam \divisor_inst.counter_0_LC_14_18_5 .C_ON=1'b0;
    defparam \divisor_inst.counter_0_LC_14_18_5 .SEQ_MODE=4'b1010;
    defparam \divisor_inst.counter_0_LC_14_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \divisor_inst.counter_0_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11996),
            .lcout(divisor_inst_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10836),
            .ce(),
            .sr(N__10628));
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_fast_1_LC_14_19_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_fast_1_LC_14_19_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_fast_1_LC_14_19_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_fast_fast_1_LC_14_19_1  (
            .in0(N__11624),
            .in1(N__11369),
            .in2(N__8498),
            .in3(N__11689),
            .lcout(\FSM_TEST_inst_RAPIDA.current_state_fast_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10845),
            .ce(),
            .sr(N__10623));
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_LC_14_19_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_LC_14_19_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_LC_14_19_2 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_fast_1_rep1_LC_14_19_2  (
            .in0(N__11366),
            .in1(N__8450),
            .in2(N__11690),
            .in3(N__11623),
            .lcout(\FSM_TEST_inst_RAPIDA.current_state_fast_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10845),
            .ce(),
            .sr(N__10623));
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_1_LC_14_19_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_1_LC_14_19_3 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_1_LC_14_19_3 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_fast_1_LC_14_19_3  (
            .in0(N__11622),
            .in1(N__11685),
            .in2(N__9411),
            .in3(N__11368),
            .lcout(\FSM_TEST_inst_RAPIDA.current_state_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10845),
            .ce(),
            .sr(N__10623));
    defparam \FSM_TEST_inst_slow.CLK_uC_6l_0_LC_14_19_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_slow.CLK_uC_6l_0_LC_14_19_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_slow.CLK_uC_6l_0_LC_14_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FSM_TEST_inst_slow.CLK_uC_6l_0_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9356),
            .lcout(CLK_uC_6l_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10845),
            .ce(),
            .sr(N__10623));
    defparam \FSM_TEST_inst_RAPIDA.current_state_1_rep1_LC_14_19_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_1_rep1_LC_14_19_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.current_state_1_rep1_LC_14_19_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_1_rep1_LC_14_19_5  (
            .in0(N__11621),
            .in1(N__11684),
            .in2(N__10243),
            .in3(N__11367),
            .lcout(\FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10845),
            .ce(),
            .sr(N__10623));
    defparam \FSM_TEST_inst_RAPIDA.counter_din_0_LC_14_19_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_din_0_LC_14_19_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.counter_din_0_LC_14_19_7 .LUT_INIT=16'b0110011001000100;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_din_0_LC_14_19_7  (
            .in0(N__11620),
            .in1(N__9877),
            .in2(_gnd_net_),
            .in3(N__11911),
            .lcout(\FSM_TEST_inst_RAPIDA.counter_dinZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10845),
            .ce(),
            .sr(N__10623));
    defparam \config_register_latched_dec_inst.DYNSR_3_LC_14_20_0 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNSR_3_LC_14_20_0 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNSR_3_LC_14_20_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \config_register_latched_dec_inst.DYNSR_3_LC_14_20_0  (
            .in0(N__9332),
            .in1(N__10073),
            .in2(_gnd_net_),
            .in3(N__9301),
            .lcout(\config_register_latched_dec_inst.DYNSRZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10853),
            .ce(N__9479),
            .sr(N__10617));
    defparam \config_register_latched_dec_inst.DYNSR_4_LC_14_20_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNSR_4_LC_14_20_1 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNSR_4_LC_14_20_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \config_register_latched_dec_inst.DYNSR_4_LC_14_20_1  (
            .in0(N__9323),
            .in1(N__10069),
            .in2(_gnd_net_),
            .in3(N__9331),
            .lcout(\config_register_latched_dec_inst.DYNSRZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10853),
            .ce(N__9479),
            .sr(N__10617));
    defparam \config_register_latched_dec_inst.DYNSR_5_LC_14_20_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNSR_5_LC_14_20_2 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNSR_5_LC_14_20_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \config_register_latched_dec_inst.DYNSR_5_LC_14_20_2  (
            .in0(N__10068),
            .in1(N__9554),
            .in2(_gnd_net_),
            .in3(N__9322),
            .lcout(\config_register_latched_dec_inst.DYNSRZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10853),
            .ce(N__9479),
            .sr(N__10617));
    defparam \config_register_latched_dec_inst.DYNSR_7_LC_14_20_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNSR_7_LC_14_20_3 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNSR_7_LC_14_20_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \config_register_latched_dec_inst.DYNSR_7_LC_14_20_3  (
            .in0(N__10070),
            .in1(N__9563),
            .in2(_gnd_net_),
            .in3(N__9544),
            .lcout(\config_register_latched_dec_inst.DYNSRZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10853),
            .ce(N__9479),
            .sr(N__10617));
    defparam \config_register_latched_dec_inst.DYNSR_2_LC_14_20_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNSR_2_LC_14_20_4 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNSR_2_LC_14_20_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \config_register_latched_dec_inst.DYNSR_2_LC_14_20_4  (
            .in0(N__10067),
            .in1(N__9302),
            .in2(_gnd_net_),
            .in3(N__9313),
            .lcout(\config_register_latched_dec_inst.DYNSRZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10853),
            .ce(N__9479),
            .sr(N__10617));
    defparam \config_register_latched_dec_inst.DYNSR_8_LC_14_20_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNSR_8_LC_14_20_5 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNSR_8_LC_14_20_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \config_register_latched_dec_inst.DYNSR_8_LC_14_20_5  (
            .in0(N__10071),
            .in1(N__9527),
            .in2(_gnd_net_),
            .in3(N__9562),
            .lcout(\config_register_latched_dec_inst.DYNSRZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10853),
            .ce(N__9479),
            .sr(N__10617));
    defparam \config_register_latched_dec_inst.DYNSR_6_LC_14_20_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNSR_6_LC_14_20_6 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNSR_6_LC_14_20_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \config_register_latched_dec_inst.DYNSR_6_LC_14_20_6  (
            .in0(N__9545),
            .in1(N__10074),
            .in2(_gnd_net_),
            .in3(N__9553),
            .lcout(\config_register_latched_dec_inst.DYNSRZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10853),
            .ce(N__9479),
            .sr(N__10617));
    defparam \config_register_latched_dec_inst.DYNSR_9_LC_14_20_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.DYNSR_9_LC_14_20_7 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst.DYNSR_9_LC_14_20_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \config_register_latched_dec_inst.DYNSR_9_LC_14_20_7  (
            .in0(N__10072),
            .in1(N__9498),
            .in2(_gnd_net_),
            .in3(N__9528),
            .lcout(\config_register_latched_dec_inst.DYNSRZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10853),
            .ce(N__9479),
            .sr(N__10617));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_31_LC_14_21_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_31_LC_14_21_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_31_LC_14_21_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_31_LC_14_21_0  (
            .in0(N__9626),
            .in1(N__11847),
            .in2(_gnd_net_),
            .in3(N__11463),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10860),
            .ce(N__12147),
            .sr(N__10613));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_52_LC_14_21_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_52_LC_14_21_1 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_52_LC_14_21_1 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_52_LC_14_21_1  (
            .in0(N__11462),
            .in1(N__11030),
            .in2(_gnd_net_),
            .in3(N__9455),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10860),
            .ce(N__12147),
            .sr(N__10613));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_51_LC_14_21_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_51_LC_14_21_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_51_LC_14_21_2 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_51_LC_14_21_2  (
            .in0(N__11461),
            .in1(N__9431),
            .in2(_gnd_net_),
            .in3(N__11851),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10860),
            .ce(N__12147),
            .sr(N__10613));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_53_LC_14_21_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_53_LC_14_21_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_53_LC_14_21_4 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_53_LC_14_21_4  (
            .in0(N__11031),
            .in1(N__9449),
            .in2(_gnd_net_),
            .in3(N__11465),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10860),
            .ce(N__12147),
            .sr(N__10613));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_32_LC_14_21_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_32_LC_14_21_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_32_LC_14_21_5 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_32_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(N__11460),
            .in2(N__11870),
            .in3(N__9437),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10860),
            .ce(N__12147),
            .sr(N__10613));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_50_LC_14_21_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_50_LC_14_21_6 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_50_LC_14_21_6 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_50_LC_14_21_6  (
            .in0(N__11029),
            .in1(N__9809),
            .in2(_gnd_net_),
            .in3(N__11464),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10860),
            .ce(N__12147),
            .sr(N__10613));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_9_LC_14_22_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_9_LC_14_22_0 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_9_LC_14_22_0 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_9_LC_14_22_0  (
            .in0(N__11469),
            .in1(N__11869),
            .in2(_gnd_net_),
            .in3(N__9593),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10867),
            .ce(N__12143),
            .sr(N__10609));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_30_LC_14_22_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_30_LC_14_22_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_30_LC_14_22_1 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_30_LC_14_22_1  (
            .in0(N__11865),
            .in1(N__9632),
            .in2(_gnd_net_),
            .in3(N__11471),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10867),
            .ce(N__12143),
            .sr(N__10609));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_75_LC_14_22_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_75_LC_14_22_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_75_LC_14_22_3 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_75_LC_14_22_3  (
            .in0(N__11033),
            .in1(N__9785),
            .in2(_gnd_net_),
            .in3(N__11473),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10867),
            .ce(N__12143),
            .sr(N__10609));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_61_LC_14_22_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_61_LC_14_22_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_61_LC_14_22_4 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_61_LC_14_22_4  (
            .in0(N__11467),
            .in1(N__11867),
            .in2(_gnd_net_),
            .in3(N__9614),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10867),
            .ce(N__12143),
            .sr(N__10609));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_58_LC_14_22_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_58_LC_14_22_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_58_LC_14_22_5 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_58_LC_14_22_5  (
            .in0(N__11866),
            .in1(N__9581),
            .in2(_gnd_net_),
            .in3(N__11472),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10867),
            .ce(N__12143),
            .sr(N__10609));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_8_LC_14_22_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_8_LC_14_22_6 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_8_LC_14_22_6 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_8_LC_14_22_6  (
            .in0(N__11468),
            .in1(N__11868),
            .in2(_gnd_net_),
            .in3(N__9602),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10867),
            .ce(N__12143),
            .sr(N__10609));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_10_LC_14_22_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_10_LC_14_22_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_10_LC_14_22_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_10_LC_14_22_7  (
            .in0(N__10244),
            .in1(N__9587),
            .in2(_gnd_net_),
            .in3(N__11470),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10867),
            .ce(N__12143),
            .sr(N__10609));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_57_LC_14_23_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_57_LC_14_23_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_57_LC_14_23_0 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_57_LC_14_23_0  (
            .in0(N__11474),
            .in1(N__11872),
            .in2(_gnd_net_),
            .in3(N__9683),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10873),
            .ce(N__12140),
            .sr(N__10605));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_80_LC_14_23_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_80_LC_14_23_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_80_LC_14_23_4 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_80_LC_14_23_4  (
            .in0(N__11475),
            .in1(N__11873),
            .in2(_gnd_net_),
            .in3(N__9575),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10873),
            .ce(N__12140),
            .sr(N__10605));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_56_LC_14_23_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_56_LC_14_23_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_56_LC_14_23_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_56_LC_14_23_7  (
            .in0(N__11871),
            .in1(N__9689),
            .in2(_gnd_net_),
            .in3(N__11476),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10873),
            .ce(N__12140),
            .sr(N__10605));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_83_LC_15_19_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_83_LC_15_19_0 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_83_LC_15_19_0 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_83_LC_15_19_0  (
            .in0(N__10968),
            .in1(N__9638),
            .in2(_gnd_net_),
            .in3(N__11456),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10837),
            .ce(N__12150),
            .sr(N__10618));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_84_LC_15_19_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_84_LC_15_19_1 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_84_LC_15_19_1 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_84_LC_15_19_1  (
            .in0(N__11454),
            .in1(N__10969),
            .in2(_gnd_net_),
            .in3(N__9677),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10837),
            .ce(N__12150),
            .sr(N__10618));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_87_LC_15_19_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_87_LC_15_19_2 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_87_LC_15_19_2 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_87_LC_15_19_2  (
            .in0(N__10972),
            .in1(N__9644),
            .in2(_gnd_net_),
            .in3(N__11458),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10837),
            .ce(N__12150),
            .sr(N__10618));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_85_LC_15_19_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_85_LC_15_19_4 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_85_LC_15_19_4 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_85_LC_15_19_4  (
            .in0(N__10970),
            .in1(N__9656),
            .in2(_gnd_net_),
            .in3(N__11457),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10837),
            .ce(N__12150),
            .sr(N__10618));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_86_LC_15_19_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_86_LC_15_19_7 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_86_LC_15_19_7 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_86_LC_15_19_7  (
            .in0(N__11455),
            .in1(N__10971),
            .in2(_gnd_net_),
            .in3(N__9650),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10837),
            .ce(N__12150),
            .sr(N__10618));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_46_LC_15_20_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_46_LC_15_20_0 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_46_LC_15_20_0 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_46_LC_15_20_0  (
            .in0(N__11496),
            .in1(N__11023),
            .in2(_gnd_net_),
            .in3(N__9833),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10846),
            .ce(N__12148),
            .sr(N__10614));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_35_LC_15_20_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_35_LC_15_20_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_35_LC_15_20_1 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_35_LC_15_20_1  (
            .in0(N__11810),
            .in1(N__9797),
            .in2(_gnd_net_),
            .in3(N__11498),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10846),
            .ce(N__12148),
            .sr(N__10614));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_82_LC_15_20_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_82_LC_15_20_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_82_LC_15_20_3 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_82_LC_15_20_3  (
            .in0(N__11025),
            .in1(N__9725),
            .in2(_gnd_net_),
            .in3(N__11501),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10846),
            .ce(N__12148),
            .sr(N__10614));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_66_LC_15_20_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_66_LC_15_20_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_66_LC_15_20_4 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_66_LC_15_20_4  (
            .in0(N__11497),
            .in1(N__11812),
            .in2(_gnd_net_),
            .in3(N__9746),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10846),
            .ce(N__12148),
            .sr(N__10614));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_65_LC_15_20_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_65_LC_15_20_5 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_65_LC_15_20_5 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_65_LC_15_20_5  (
            .in0(N__11024),
            .in1(N__10406),
            .in2(_gnd_net_),
            .in3(N__11500),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10846),
            .ce(N__12148),
            .sr(N__10614));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_36_LC_15_20_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_36_LC_15_20_6 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_36_LC_15_20_6 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_36_LC_15_20_6  (
            .in0(N__11495),
            .in1(N__11022),
            .in2(_gnd_net_),
            .in3(N__9740),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10846),
            .ce(N__12148),
            .sr(N__10614));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_40_LC_15_20_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_40_LC_15_20_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_40_LC_15_20_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_40_LC_15_20_7  (
            .in0(N__11811),
            .in1(N__9713),
            .in2(_gnd_net_),
            .in3(N__11499),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10846),
            .ce(N__12148),
            .sr(N__10614));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_81_LC_15_21_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_81_LC_15_21_0 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_81_LC_15_21_0 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_81_LC_15_21_0  (
            .in0(N__11505),
            .in1(N__11028),
            .in2(_gnd_net_),
            .in3(N__9734),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10854),
            .ce(N__12144),
            .sr(N__10610));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_33_LC_15_21_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_33_LC_15_21_1 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_33_LC_15_21_1 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_33_LC_15_21_1  (
            .in0(N__11026),
            .in1(N__9719),
            .in2(_gnd_net_),
            .in3(N__11506),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10854),
            .ce(N__12144),
            .sr(N__10610));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_39_LC_15_21_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_39_LC_15_21_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_39_LC_15_21_2 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_39_LC_15_21_2  (
            .in0(N__11502),
            .in1(N__11832),
            .in2(_gnd_net_),
            .in3(N__9827),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10854),
            .ce(N__12144),
            .sr(N__10610));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_48_LC_15_21_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_48_LC_15_21_3 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_48_LC_15_21_3 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_48_LC_15_21_3  (
            .in0(N__11835),
            .in1(N__9701),
            .in2(_gnd_net_),
            .in3(N__11509),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10854),
            .ce(N__12144),
            .sr(N__10610));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_47_LC_15_21_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_47_LC_15_21_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_47_LC_15_21_4 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_47_LC_15_21_4  (
            .in0(N__11503),
            .in1(N__11834),
            .in2(_gnd_net_),
            .in3(N__9707),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10854),
            .ce(N__12144),
            .sr(N__10610));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_41_LC_15_21_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_41_LC_15_21_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_41_LC_15_21_5 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_41_LC_15_21_5  (
            .in0(N__11833),
            .in1(N__9695),
            .in2(_gnd_net_),
            .in3(N__11508),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10854),
            .ce(N__12144),
            .sr(N__10610));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_49_LC_15_21_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_49_LC_15_21_6 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_49_LC_15_21_6 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_49_LC_15_21_6  (
            .in0(N__11504),
            .in1(N__11027),
            .in2(_gnd_net_),
            .in3(N__9815),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10854),
            .ce(N__12144),
            .sr(N__10610));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_34_LC_15_21_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_34_LC_15_21_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_34_LC_15_21_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_34_LC_15_21_7  (
            .in0(N__11831),
            .in1(N__9803),
            .in2(_gnd_net_),
            .in3(N__11507),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10854),
            .ce(N__12144),
            .sr(N__10610));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_11_LC_15_22_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_11_LC_15_22_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_11_LC_15_22_0 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_11_LC_15_22_0  (
            .in0(N__11513),
            .in1(N__10306),
            .in2(_gnd_net_),
            .in3(N__9791),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10861),
            .ce(N__12141),
            .sr(N__10606));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_74_LC_15_22_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_74_LC_15_22_1 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_74_LC_15_22_1 .LUT_INIT=16'b1110111010111011;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_74_LC_15_22_1  (
            .in0(N__12158),
            .in1(N__11032),
            .in2(_gnd_net_),
            .in3(N__11520),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10861),
            .ce(N__12141),
            .sr(N__10606));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_16_LC_15_22_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_16_LC_15_22_2 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_16_LC_15_22_2 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_16_LC_15_22_2  (
            .in0(N__11515),
            .in1(N__11853),
            .in2(_gnd_net_),
            .in3(N__9767),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10861),
            .ce(N__12141),
            .sr(N__10606));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_13_LC_15_22_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_13_LC_15_22_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_13_LC_15_22_3 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_13_LC_15_22_3  (
            .in0(N__11852),
            .in1(N__10163),
            .in2(_gnd_net_),
            .in3(N__11518),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10861),
            .ce(N__12141),
            .sr(N__10606));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_14_LC_15_22_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_14_LC_15_22_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_14_LC_15_22_4 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_14_LC_15_22_4  (
            .in0(N__11514),
            .in1(N__10308),
            .in2(_gnd_net_),
            .in3(N__9779),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10861),
            .ce(N__12141),
            .sr(N__10606));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_15_LC_15_22_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_15_LC_15_22_5 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_15_LC_15_22_5 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_15_LC_15_22_5  (
            .in0(N__10309),
            .in1(N__9773),
            .in2(_gnd_net_),
            .in3(N__11519),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10861),
            .ce(N__12141),
            .sr(N__10606));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_17_LC_15_22_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_17_LC_15_22_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_17_LC_15_22_6 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_17_LC_15_22_6  (
            .in0(N__11516),
            .in1(N__10310),
            .in2(_gnd_net_),
            .in3(N__9761),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10861),
            .ce(N__12141),
            .sr(N__10606));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_12_LC_15_22_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_12_LC_15_22_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_12_LC_15_22_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_12_LC_15_22_7  (
            .in0(N__10307),
            .in1(N__10169),
            .in2(_gnd_net_),
            .in3(N__11517),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10861),
            .ce(N__12141),
            .sr(N__10606));
    defparam \config_register_latched_dec_inst.STATCNF_1_RNIRDN51_0_LC_16_19_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.STATCNF_1_RNIRDN51_0_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst.STATCNF_1_RNIRDN51_0_LC_16_19_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \config_register_latched_dec_inst.STATCNF_1_RNIRDN51_0_LC_16_19_1  (
            .in0(N__12097),
            .in1(N__10157),
            .in2(N__10130),
            .in3(N__10094),
            .lcout(\config_register_latched_dec_inst.STATCNF_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.counter_din_RNIEMB2_3_LC_16_19_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.counter_din_RNIEMB2_3_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.counter_din_RNIEMB2_3_LC_16_19_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.counter_din_RNIEMB2_3_LC_16_19_3  (
            .in0(N__9972),
            .in1(N__9941),
            .in2(N__9911),
            .in3(N__9881),
            .lcout(\FSM_TEST_inst_RAPIDA.N_123_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_68_LC_16_20_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_68_LC_16_20_0 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_68_LC_16_20_0 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_68_LC_16_20_0  (
            .in0(N__10944),
            .in1(N__9839),
            .in2(_gnd_net_),
            .in3(N__11512),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10831),
            .ce(N__12145),
            .sr(N__10607));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_67_LC_16_20_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_67_LC_16_20_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_67_LC_16_20_3 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_67_LC_16_20_3  (
            .in0(N__11510),
            .in1(N__10943),
            .in2(_gnd_net_),
            .in3(N__9845),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10831),
            .ce(N__12145),
            .sr(N__10607));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_45_LC_16_20_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_45_LC_16_20_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_45_LC_16_20_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_45_LC_16_20_6  (
            .in0(N__11723),
            .in1(N__10412),
            .in2(_gnd_net_),
            .in3(N__11511),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10831),
            .ce(N__12145),
            .sr(N__10607));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_38_LC_16_21_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_38_LC_16_21_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_38_LC_16_21_0 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_38_LC_16_21_0  (
            .in0(N__11521),
            .in1(N__11824),
            .in2(_gnd_net_),
            .in3(N__10424),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10840),
            .ce(N__12142),
            .sr(N__10604));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_43_LC_16_21_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_43_LC_16_21_2 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_43_LC_16_21_2 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_43_LC_16_21_2  (
            .in0(N__11522),
            .in1(_gnd_net_),
            .in2(N__10364),
            .in3(N__11825),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10840),
            .ce(N__12142),
            .sr(N__10604));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_37_LC_16_21_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_37_LC_16_21_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_37_LC_16_21_3 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_37_LC_16_21_3  (
            .in0(N__10999),
            .in1(N__9821),
            .in2(_gnd_net_),
            .in3(N__11524),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10840),
            .ce(N__12142),
            .sr(N__10604));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_44_LC_16_21_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_44_LC_16_21_5 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_44_LC_16_21_5 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_44_LC_16_21_5  (
            .in0(N__11000),
            .in1(N__10418),
            .in2(_gnd_net_),
            .in3(N__11525),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10840),
            .ce(N__12142),
            .sr(N__10604));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_64_LC_16_21_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_64_LC_16_21_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_64_LC_16_21_6 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_64_LC_16_21_6  (
            .in0(N__11523),
            .in1(N__11826),
            .in2(_gnd_net_),
            .in3(N__10400),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10840),
            .ce(N__12142),
            .sr(N__10604));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_63_LC_16_21_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_63_LC_16_21_7 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_63_LC_16_21_7 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_63_LC_16_21_7  (
            .in0(N__11001),
            .in1(N__10385),
            .in2(_gnd_net_),
            .in3(N__11526),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10840),
            .ce(N__12142),
            .sr(N__10604));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_62_LC_16_22_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_62_LC_16_22_1 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_62_LC_16_22_1 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_62_LC_16_22_1  (
            .in0(N__11827),
            .in1(N__10394),
            .in2(_gnd_net_),
            .in3(N__11531),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10848),
            .ce(N__12139),
            .sr(N__10603));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_69_LC_16_22_2 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_69_LC_16_22_2 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_69_LC_16_22_2 .LUT_INIT=16'b1111111110011001;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_69_LC_16_22_2  (
            .in0(N__11527),
            .in1(N__11003),
            .in2(_gnd_net_),
            .in3(N__10379),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10848),
            .ce(N__12139),
            .sr(N__10603));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_42_LC_16_22_3 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_42_LC_16_22_3 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_42_LC_16_22_3 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_42_LC_16_22_3  (
            .in0(N__11002),
            .in1(N__10370),
            .in2(_gnd_net_),
            .in3(N__11530),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10848),
            .ce(N__12139),
            .sr(N__10603));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_70_LC_16_22_4 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_70_LC_16_22_4 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_70_LC_16_22_4 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_70_LC_16_22_4  (
            .in0(N__11528),
            .in1(N__11828),
            .in2(_gnd_net_),
            .in3(N__10355),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10848),
            .ce(N__12139),
            .sr(N__10603));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_71_LC_16_22_5 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_71_LC_16_22_5 .SEQ_MODE=4'b1011;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_71_LC_16_22_5 .LUT_INIT=16'b1110111011011101;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_71_LC_16_22_5  (
            .in0(N__11004),
            .in1(N__10349),
            .in2(_gnd_net_),
            .in3(N__11532),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10848),
            .ce(N__12139),
            .sr(N__10603));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_72_LC_16_22_6 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_72_LC_16_22_6 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_72_LC_16_22_6 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_72_LC_16_22_6  (
            .in0(N__11529),
            .in1(N__11829),
            .in2(_gnd_net_),
            .in3(N__12170),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10848),
            .ce(N__12139),
            .sr(N__10603));
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_73_LC_16_22_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_73_LC_16_22_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.bit_sequence_stat_73_LC_16_22_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.bit_sequence_stat_73_LC_16_22_7  (
            .in0(N__11830),
            .in1(N__12164),
            .in2(_gnd_net_),
            .in3(N__11533),
            .lcout(\FSM_TEST_inst_RAPIDA.bit_sequence_statZ0Z_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10848),
            .ce(N__12139),
            .sr(N__10603));
    defparam RST_N_ibuf_RNIBJGC_LC_16_30_0.C_ON=1'b0;
    defparam RST_N_ibuf_RNIBJGC_LC_16_30_0.SEQ_MODE=4'b0000;
    defparam RST_N_ibuf_RNIBJGC_LC_16_30_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 RST_N_ibuf_RNIBJGC_LC_16_30_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12034),
            .lcout(RST_N_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIKIU51_1_LC_17_18_1 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIKIU51_1_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIKIU51_1_LC_17_18_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIKIU51_1_LC_17_18_1  (
            .in0(N__11999),
            .in1(N__11968),
            .in2(N__11939),
            .in3(N__11912),
            .lcout(\FSM_TEST_inst_RAPIDA.current_state_fast_fast_RNIKIU51Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FSM_TEST_inst_RAPIDA.current_state_1_rep2_LC_17_19_0 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_1_rep2_LC_17_19_0 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.current_state_1_rep2_LC_17_19_0 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_1_rep2_LC_17_19_0  (
            .in0(N__11493),
            .in1(N__11671),
            .in2(N__11749),
            .in3(N__11656),
            .lcout(\FSM_TEST_inst_RAPIDA.current_state_1_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10838),
            .ce(),
            .sr(N__10619));
    defparam \FSM_TEST_inst_RAPIDA.current_state_1_LC_17_19_7 .C_ON=1'b0;
    defparam \FSM_TEST_inst_RAPIDA.current_state_1_LC_17_19_7 .SEQ_MODE=4'b1010;
    defparam \FSM_TEST_inst_RAPIDA.current_state_1_LC_17_19_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \FSM_TEST_inst_RAPIDA.current_state_1_LC_17_19_7  (
            .in0(N__11670),
            .in1(N__11655),
            .in2(N__10967),
            .in3(N__11494),
            .lcout(\FSM_TEST_inst_RAPIDA.current_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10838),
            .ce(),
            .sr(N__10619));
    defparam \config_register_latched_dec_inst.STATCNF_1_RNIRDN51_0_0_LC_20_19_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst.STATCNF_1_RNIRDN51_0_0_LC_20_19_1 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst.STATCNF_1_RNIRDN51_0_0_LC_20_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \config_register_latched_dec_inst.STATCNF_1_RNIRDN51_0_0_LC_20_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10454),
            .lcout(STATCNF_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
