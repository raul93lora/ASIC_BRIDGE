/* 
* Raul Lora Rivera
* Module that send the DYNCNF and STATCNF to analog part of ASIC at 1MHz frequency
*
*/
module switch_clk_1MHz #(
    parameter DELAY_CYCLES = 17,
    parameter BIT_SEQUENCE_DIN_INIT = 16'hABC6,   				// DYNCNF default value
    parameter BIT_SEQUENCE_STAT_INIT = 88'h123456789ABCDEF1234567  	// STATCNF default value
)(
	CLK,									// Faster clock: f_CLK > f_clk_continuous_1MHz
	clk_continuous_1MHz,							// Continuous clk (1MHz), slower than CLK
	CLK_ON_OFF,								// ON/OFF clock (activated/deactivated in the corresponding states)
	RST_N,									// Low active reset
	SEL,									// Signal to choose between dynamic or static register
	flag_input,
	MOSI 									// Master Output - Slave Input
);

	// Size parameters definition
	parameter SIZESRSTAT = 88; 						// Static shift register length 
	parameter SIZESRDYN = 16; 						// Dynamic shift register length

	// Wait parameters definition
	parameter N_CYCLES_IDLE = 200; 					// Clock cycles to wait in IDLE
	parameter N_CYCLES_DYN_READ = 16; 					// Dynamic register length WAIT
	parameter N_CYCLES_STATIC_READ = 88;					// Static register length WAIT

    	// Ports definition
	input wire flag_input;
	reg flag_input_reg;
    	input wire CLK;
	input wire clk_continuous_1MHz;
	input wire RST_N;
	output reg SEL;
	output reg MOSI;
	output wire CLK_ON_OFF;
	
	// Reg signals
	reg CLK_uC;

    	// Parameters definition -- Definition of states
    	parameter IDLE = 3'b000;
    	parameter DYN_READ = 3'b001;
    	parameter STATIC_READ = 3'b010;
	parameter INDEF_STATE = 3'b011;

    	// Waiting counters in IDLE, DYN_READ y STATIC_READ states
    	reg [13:0] counter_idle; 						// 10-bit counter (up to 1024 cycles)
    	reg [3:0] counter_din;						// 4-bit counter (up to 16 cycles)
    	reg [6:0] counter_stat;						// 7-bit counter (up to 128 cycles), although only 89 are needed

    	// Current and next states
    	reg [2:0] current_state, next_state;

    	// Registers to store the dynamic and static bit sequences
    	reg [15:0] bit_sequence_din;  					// Store 16 bits for dynamic register
	reg [87:0] bit_sequence_stat;	  					// Store 89 bits for static register

	// Sequential assignment of aux_CLK
	always @(posedge CLK or negedge RST_N) begin
		if(!RST_N) begin
			CLK_uC <= 0;
		end else if (current_state == DYN_READ || current_state == STATIC_READ) begin
			CLK_uC <= clk_continuous_1MHz;
		end
	end	

	// Delay of 17 CLK cycles to ahieve the 1MHz frequency
	delay_chain #(
    		.DELAY_CYCLES(DELAY_CYCLES)
	) delay_inst (
    		.clk(CLK),
    		.rst_n(RST_N),
    		.in_signal(CLK_uC),
    		.out_signal(CLK_ON_OFF)
	);

	// Sequential assignment for flag_input signal
	always @(posedge CLK or negedge RST_N) begin
		if(!RST_N) begin
			flag_input_reg <= 0;
		end else begin
			flag_input_reg <= flag_input;
		end
	end

    	// State-transition logic
    	always @(posedge clk_continuous_1MHz or negedge RST_N) begin
        	if (!RST_N) begin
            		current_state <= IDLE; 				// When reset, it goes to IDLE state
        	end else begin
            		current_state <= next_state; 				// Next state change
        	end
    	end

    	// Next State logic
    	always @(*) begin
        	case (current_state)
            		IDLE: next_state = (flag_input_reg == 1 && counter_idle >= N_CYCLES_IDLE-1) ? DYN_READ : IDLE;			// From IDLE, it goes to DYN_READ, after waiting for N_CYCLES_IDLE
            		DYN_READ: next_state = (counter_din == N_CYCLES_DYN_READ-1) ? STATIC_READ : DYN_READ;				// From DYN_READ, it goes to STATIC_READ, after waiting for N_CYCLES_DYN_READ
            		STATIC_READ: next_state = (counter_stat == N_CYCLES_STATIC_READ-1) ? INDEF_STATE : STATIC_READ;		// From STATIC_READ, it goes to INDEF_STATE, after waiting for N_CYCLES_STATIC_READ
			INDEF_STATE: next_state = INDEF_STATE;										// It has to wait indefinitely in order to have the correct behaviour
            		default: next_state = IDLE;												// Default: Vuelve a IDLE
        	endcase
    	end

	// Output logic - FSM
	always @(posedge clk_continuous_1MHz or negedge RST_N) begin
		if (!RST_N) begin
			SEL <= 0;
			MOSI <= 0;
			bit_sequence_din <= BIT_SEQUENCE_DIN_INIT; 
			bit_sequence_stat <= BIT_SEQUENCE_STAT_INIT;			
		end else begin
            	case (current_state)
			IDLE: begin
				SEL <= 0;
				MOSI <= 0;
				bit_sequence_din <= BIT_SEQUENCE_DIN_INIT; 
				bit_sequence_stat <= BIT_SEQUENCE_STAT_INIT;
			end
			DYN_READ: begin
				SEL <= 1;	
                    		// Shift sequence and update output signal
                    		MOSI <= bit_sequence_din[SIZESRDYN-1]; 					// El bit m�s significativo de la secuencia
                    		bit_sequence_din <= {bit_sequence_din[SIZESRDYN-2:0], 1'b0};  	// Desplazamos la secuencia a la izquierda
               	end
               	STATIC_READ: begin
				SEL <= 0;
                    		// Shift sequence and update output signal
                    		MOSI <= bit_sequence_stat[SIZESRSTAT-1]; 					// The most significant bit of the sequence								
                    		bit_sequence_stat <= {bit_sequence_stat[SIZESRSTAT-2:0], 1'b0};  		// Left-Shift the sequence
               	end
			INDEF_STATE: begin									// It has to wait indefinitely in this state
				SEL <= 1;
				MOSI <= 0;
				bit_sequence_din <= BIT_SEQUENCE_DIN_INIT; 
				bit_sequence_stat <= BIT_SEQUENCE_STAT_INIT;
			end
               	default: begin
				SEL <= 0;
				MOSI <= 0;
				bit_sequence_din <= BIT_SEQUENCE_DIN_INIT; 
				bit_sequence_stat <= BIT_SEQUENCE_STAT_INIT;
               	end
            	endcase
        	end
    	end

    	// Counter to wait in IDLE state
    	always @(posedge clk_continuous_1MHz or negedge RST_N) begin
       		if (!RST_N) begin
            		counter_idle <= 0; 							  		// Reset the counter
        	end else if (current_state == IDLE && counter_idle < N_CYCLES_IDLE) begin
            		counter_idle <= counter_idle + 1; 							// Increase the counter in IDLE state
        	end else if (current_state != IDLE) begin
            		counter_idle <= 0; 									// Reset counter when no IDLE state
        	end
    	end

    	// Counter to wait in DYN_READ state
    	always @(posedge clk_continuous_1MHz or negedge RST_N) begin
       		if (!RST_N) begin
            		counter_din <= 0; 							  		// Reset the counter
        	end else if (current_state == DYN_READ && counter_din < N_CYCLES_DYN_READ) begin
            		counter_din <= counter_din + 1; 							// Increase the counter in DYN_READ state
        	end else if (current_state != DYN_READ) begin
            		counter_din <= 0; 									// Reset counter when no DYN_READ state
        	end
    	end

    	// Counter to wait in STATIC_READ state
    	always @(posedge clk_continuous_1MHz or negedge RST_N) begin
       		if (!RST_N) begin
            		counter_stat <= 0; 							  		// Reset the counter
        	end else if (current_state == STATIC_READ && counter_stat < N_CYCLES_STATIC_READ) begin
            		counter_stat <= counter_stat + 1; 							// Increase the counter in STATIC_READ
        	end else if (current_state != STATIC_READ) begin
            		counter_stat <= 0; 									// Reset counter when no STATIC_READ state
        	end
    	end   

endmodule








