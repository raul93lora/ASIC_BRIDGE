-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     May 15 2025 16:30:08

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "ASIC_bridge_top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of ASIC_bridge_top
entity ASIC_bridge_top is
port (
    xor_out_dyn : out std_logic;
    sel_output : out std_logic;
    clk_output : out std_logic;
    CLK : in std_logic;
    xor_out_stat : out std_logic;
    mosi_output : out std_logic;
    miso_input : in std_logic;
    RST_N : in std_logic);
end ASIC_bridge_top;

-- Architecture of ASIC_bridge_top
-- View name is \INTERFACE\
architecture \INTERFACE\ of ASIC_bridge_top is

signal \N__11095\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \CLK_ibuf_gb_io_gb_input\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_13\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_12\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_79\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_11\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_78\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_10\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_55\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_76\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_77\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_36\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_53\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_54\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_5\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_6\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_7\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_8\ : std_logic;
signal \RST_N_c_i\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_14\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_15\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_73\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_9\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_56\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_57\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_27\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_44\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_26\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_35\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_34\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_37\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_43\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_52\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_74\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_75\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_16\ : std_logic;
signal \switch_clk_2MHz_inst.counter_idlelde_2_cascade_\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_0\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_1\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_2\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_3\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_4\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_13\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_14\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_12\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_9\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_10\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_11\ : std_logic;
signal \switch_clk_2MHz_inst.current_state_fast_RNIJRTPZ0Z_1\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_6\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_2\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_7\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_0\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_1\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_3\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_4\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_5\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_68\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_80\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_64\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_65\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_8\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_21\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_66\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_67\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_30\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_28\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_29\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_38\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_20\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_19\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_33\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_31\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_32\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_42\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_17\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_18\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_50\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_51\ : std_logic;
signal \switch_clk_2MHz_inst.aux_CLKZ0\ : std_logic;
signal \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_0\ : std_logic;
signal \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_1\ : std_logic;
signal \bfn_3_21_0_\ : std_logic;
signal \switch_clk_2MHz_inst.counter_idle_cry_0\ : std_logic;
signal \switch_clk_2MHz_inst.counter_idle_cry_1\ : std_logic;
signal \switch_clk_2MHz_inst.counter_idle_cry_2\ : std_logic;
signal \switch_clk_2MHz_inst.counter_idle_cry_3\ : std_logic;
signal \switch_clk_2MHz_inst.counter_idle_cry_4\ : std_logic;
signal \switch_clk_2MHz_inst.current_state_fast_RNIDHKD1Z0Z_1\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_8\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_9\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_10\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_11\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_14\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_12\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_13\ : std_logic;
signal \switch_clk_1MHz_inst.counter_statlde_0_cascade_\ : std_logic;
signal \switch_clk_1MHz_inst.current_state_RNITOE91Z0Z_1\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_72\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_81\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_69\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_70\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_71\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_22\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_62\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_63\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_58\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_23\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_4\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_49\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_45\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_7\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_24\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_25\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_3\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_0\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_1\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_2\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_5\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_6\ : std_logic;
signal \switch_clk_2MHz_inst.counter_statZ0Z_0\ : std_logic;
signal \bfn_4_20_0_\ : std_logic;
signal \switch_clk_2MHz_inst.counter_stat_cry_0\ : std_logic;
signal \switch_clk_2MHz_inst.counter_statZ0Z_2\ : std_logic;
signal \switch_clk_2MHz_inst.counter_stat_cry_1\ : std_logic;
signal \switch_clk_2MHz_inst.counter_stat_cry_2\ : std_logic;
signal \switch_clk_2MHz_inst.counter_stat_cry_3\ : std_logic;
signal \switch_clk_2MHz_inst.counter_stat_cry_4\ : std_logic;
signal \switch_clk_2MHz_inst.counter_stat_cry_5\ : std_logic;
signal \switch_clk_2MHz_inst.counter_idleZ0Z_0\ : std_logic;
signal \switch_clk_2MHz_inst.counter_idleZ0Z_1\ : std_logic;
signal \switch_clk_2MHz_inst.counter_idleZ0Z_2\ : std_logic;
signal \switch_clk_2MHz_inst.counter_idleZ0Z_5\ : std_logic;
signal \switch_clk_2MHz_inst.counter_idleZ0Z_4\ : std_logic;
signal \switch_clk_2MHz_inst.counter_idleZ0Z_3\ : std_logic;
signal \switch_clk_2MHz_inst.G_31_0_a4_0_4\ : std_logic;
signal \switch_clk_2MHz_inst.G_31_0_a4_0_5_cascade_\ : std_logic;
signal \switch_clk_1MHz_inst.current_state_ns_0_a3_1_4_0_cascade_\ : std_logic;
signal \switch_clk_2MHz_inst.N_117_1_i\ : std_logic;
signal \switch_clk_1MHz_inst.counter_statZ0Z_0\ : std_logic;
signal \bfn_4_22_0_\ : std_logic;
signal \switch_clk_1MHz_inst.counter_stat_cry_0\ : std_logic;
signal \switch_clk_1MHz_inst.counter_statZ0Z_2\ : std_logic;
signal \switch_clk_1MHz_inst.counter_stat_cry_1\ : std_logic;
signal \switch_clk_1MHz_inst.counter_statZ0Z_3\ : std_logic;
signal \switch_clk_1MHz_inst.counter_stat_cry_2\ : std_logic;
signal \switch_clk_1MHz_inst.counter_stat_cry_3\ : std_logic;
signal \switch_clk_1MHz_inst.counter_stat_cry_4\ : std_logic;
signal \switch_clk_1MHz_inst.counter_stat_cry_5\ : std_logic;
signal \switch_clk_1MHz_inst.counter_statZ0Z_6\ : std_logic;
signal \switch_clk_1MHz_inst.current_state_RNIFA8B2Z0Z_1\ : std_logic;
signal \bfn_4_23_0_\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idle_cry_0\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idle_cry_1\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idle_cry_2\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idle_cry_3\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idle_cry_4\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idle_cry_5\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idle_cry_6\ : std_logic;
signal \switch_clk_1MHz_inst.N_116_1\ : std_logic;
signal \switch_clk_1MHz_inst.G_31_1_cascade_\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idle_RNIOJRU1Z0Z_7\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idleZ0Z_3\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idleZ0Z_4\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idleZ0Z_7\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idleZ0Z_6\ : std_logic;
signal \switch_clk_1MHz_inst.current_state_RNO_5Z0Z_0\ : std_logic;
signal \switch_clk_1MHz_inst.current_state_RNO_4Z0Z_0_cascade_\ : std_logic;
signal \switch_clk_1MHz_inst.N_116_cascade_\ : std_logic;
signal \switch_clk_1MHz_inst.current_state_RNO_1Z0Z_0\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_58\ : std_logic;
signal \DYNCNF_i_0\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_82\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_61\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_46\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_59\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_60\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_47\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_48\ : std_logic;
signal \switch_clk_2MHz_inst.flag_input_regZ0\ : std_logic;
signal \switch_clk_2MHz_inst.N_114_0_cascade_\ : std_logic;
signal \switch_clk_2MHz_inst.current_state_1_repZ0Z1\ : std_logic;
signal \switch_clk_2MHz_inst.current_state_d_i_2\ : std_logic;
signal \switch_clk_2MHz_inst.counter_statZ0Z_3\ : std_logic;
signal \switch_clk_2MHz_inst.current_state_fastZ0Z_1\ : std_logic;
signal \switch_clk_2MHz_inst.counter_statlde_0_cascade_\ : std_logic;
signal \switch_clk_2MHz_inst.current_state_fast_RNI9DAU1Z0Z_1\ : std_logic;
signal \switch_clk_2MHz_inst.counter_statZ0Z_1\ : std_logic;
signal \switch_clk_2MHz_inst.counter_statZ0Z_6\ : std_logic;
signal \switch_clk_2MHz_inst.counter_statZ0Z_5\ : std_logic;
signal \switch_clk_2MHz_inst.counter_statZ0Z_4\ : std_logic;
signal \switch_clk_2MHz_inst.G_31_0_a4_1_1_cascade_\ : std_logic;
signal \switch_clk_2MHz_inst.G_31_0_a4_1_5\ : std_logic;
signal \switch_clk_2MHz_inst.N_9_1\ : std_logic;
signal \switch_clk_2MHz_inst.G_31_0_a4_1_6_cascade_\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idleZ0Z_2\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idleZ0Z_1\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idleZ0Z_5\ : std_logic;
signal \switch_clk_1MHz_inst.counter_idleZ0Z_0\ : std_logic;
signal \switch_clk_1MHz_inst.current_state_RNO_3Z0Z_0\ : std_logic;
signal \switch_clk_1MHz_inst.counter_statZ0Z_4\ : std_logic;
signal \switch_clk_1MHz_inst.counter_statZ0Z_1\ : std_logic;
signal \switch_clk_1MHz_inst.counter_statZ0Z_5\ : std_logic;
signal \switch_clk_1MHz_inst.current_state_ns_0_a3_1_5_0\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_15\ : std_logic;
signal \switch_clk_2MHz_inst.N_8_0\ : std_logic;
signal \switch_clk_1MHz_inst.current_state_d_i_2\ : std_logic;
signal \switch_clk_1MHz_inst.N_116_1_i\ : std_logic;
signal \config_register_latched_dec_inst.DYNCNF_0\ : std_logic;
signal \config_register_latched_dec_inst.DYNCNF_1Z0Z_0\ : std_logic;
signal \counter_RNISR1F_2_cascade_\ : std_logic;
signal \switch_clk_1MHz_inst.current_state_RNITOE91_0Z0Z_1\ : std_logic;
signal \switch_clk_1MHz_inst.current_state_cnv_0_1_cascade_\ : std_logic;
signal \switch_clk_1MHz_inst.counter_dinZ1Z_1\ : std_logic;
signal \switch_clk_1MHz_inst.counter_dinZ0Z_0\ : std_logic;
signal \switch_clk_1MHz_inst.current_state_RNO_8Z0Z_0_cascade_\ : std_logic;
signal \switch_clk_1MHz_inst.current_state_RNO_2Z0Z_0\ : std_logic;
signal \switch_clk_1MHz_inst.N_88_0\ : std_logic;
signal \switch_clk_1MHz_inst.counter_dinZ0Z_2\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_24\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_28\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_57\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_23\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_27\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_25\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_26\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_59\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_60\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_61\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_29\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_30\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_83\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_84\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_41\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_87\ : std_logic;
signal \switch_clk_2MHz_inst.current_state_1_repZ0Z2\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_39\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_40\ : std_logic;
signal \switch_clk_2MHz_inst.current_stateZ0Z_1\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_85\ : std_logic;
signal \switch_clk_2MHz_inst.bit_sequence_statZ0Z_86\ : std_logic;
signal \switch_clk_2MHz_inst.N_259_g\ : std_logic;
signal \switch_clk_2MHz_inst.counter_din_3_i_0_2_cascade_\ : std_logic;
signal \clk_out_RNI3LEM_cascade_\ : std_logic;
signal \switch_clk_2MHz_inst.G_31_0_o4_2\ : std_logic;
signal \switch_clk_2MHz_inst.counter_dinZ0Z_0\ : std_logic;
signal \switch_clk_2MHz_inst.counter_dinZ1Z_1\ : std_logic;
signal \switch_clk_2MHz_inst.counter_dinZ0Z_2\ : std_logic;
signal \switch_clk_2MHz_inst.N_92_0\ : std_logic;
signal \switch_clk_2MHz_inst.N_92_0_cascade_\ : std_logic;
signal \switch_clk_2MHz_inst.counter_dinZ0Z_3\ : std_logic;
signal \switch_clk_2MHz_inst.SEL_0_RNIC97QZ0_cascade_\ : std_logic;
signal \switch_clk_2MHz_inst.SEL_0_RNIC97QZ0Z_0\ : std_logic;
signal \switch_clk_2MHz_inst.SEL_0_RNIC97QZ0Z_0_cascade_\ : std_logic;
signal \switch_clk_2MHz_inst.SEL_0_RNIC97QZ0\ : std_logic;
signal \switch_clk_2MHz_inst.N_91_li_cascade_\ : std_logic;
signal \clk_continuous_2MHz\ : std_logic;
signal \switch_clk_2MHz_inst.current_state_fast_fast_RNI0KTVZ0Z_1\ : std_logic;
signal \switch_clk_2MHz_inst.N_114_0\ : std_logic;
signal \switch_clk_2MHz_inst.current_state_fast_fastZ0Z_1\ : std_logic;
signal \mosi_2MHz\ : std_logic;
signal mosi_output_c : std_logic;
signal \switch_clk_2MHz_inst.aux_selection_2MHz_0\ : std_logic;
signal \switch_clk_2MHz_inst.N_91_li\ : std_logic;
signal \switch_clk_2MHz_inst.SEL_0_RNI98MZ0Z31_cascade_\ : std_logic;
signal \N_381_i\ : std_logic;
signal \aux_selection_1MHz_0\ : std_logic;
signal \N_4_0_cascade_\ : std_logic;
signal \config_register_latched_dec_inst.STATCNF_1_RNO_0Z0Z_0\ : std_logic;
signal \N_2_0\ : std_logic;
signal \switch_clk_2MHz_inst.current_stateZ0Z_0\ : std_logic;
signal \switch_clk_2MHz_inst.current_state_fast_1_repZ0Z1\ : std_logic;
signal \clk_out_RNI3LEM\ : std_logic;
signal \divisor_inst_2.counterZ0Z_0\ : std_logic;
signal \divisor_inst_2.counterZ0Z_2\ : std_logic;
signal \divisor_inst_2.counterZ0Z_1\ : std_logic;
signal \switch_clk_2MHz_inst.SEL_0_RNI98MZ0Z31\ : std_logic;
signal \N_3_0\ : std_logic;
signal flag_signal : std_logic;
signal \switch_clk_1MHz_inst.flag_input_regZ0\ : std_logic;
signal \clk_continuous_1MHz\ : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_1\ : std_logic;
signal \switch_clk_1MHz_inst.N_91_0\ : std_logic;
signal \switch_clk_1MHz_inst.N_90_li\ : std_logic;
signal \switch_clk_1MHz_inst.counter_dinZ0Z_3\ : std_logic;
signal \switch_clk_1MHz_inst.CLK_uCZ0\ : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_0\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_55\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_56\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_62\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_63\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_31\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal divisor_inst_counter_1 : std_logic;
signal divisor_inst_counter_0 : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_reg_0_6\ : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_5\ : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_4\ : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_7\ : std_logic;
signal \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_2\ : std_logic;
signal \N_4_0\ : std_logic;
signal clk_output_c : std_logic;
signal \switch_clk_2MHz_inst_delay_inst_delay_reg_6\ : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_2\ : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_3\ : std_logic;
signal \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_3\ : std_logic;
signal \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_4\ : std_logic;
signal \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_5\ : std_logic;
signal \config_register_latched_dec_inst.N_381_i_i\ : std_logic;
signal \config_register_latched_dec_inst.DYNSRZ0Z_0\ : std_logic;
signal miso_input_c : std_logic;
signal \delay_reg_RNI7S8U1_15\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_32\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_54\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_12\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_13\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_14\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_52\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_53\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_11\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_9\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_10\ : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_8\ : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_9\ : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_10\ : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_11\ : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_12\ : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_13\ : std_logic;
signal \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_14\ : std_logic;
signal \switch_clk_1MHz_inst_delay_inst_delay_reg_15\ : std_logic;
signal \config_register_latched_dec_inst.STATCNF_1Z0Z_0\ : std_logic;
signal \RST_N_c\ : std_logic;
signal sel_output_c : std_logic;
signal \config_register_latched_dec_inst.STATSRZ0Z_0\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_81\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_86\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_49\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_48\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_15\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_50\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_51\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_33\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_34\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_66\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_64\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_65\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_74\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_75\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_67\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_42\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_43\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_44\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_45\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_46\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_47\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_68\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_69\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_70\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_15\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_87\ : std_logic;
signal \mosi_1MHz\ : std_logic;
signal \counter_RNISR1F_2\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_85\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_82\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_83\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_84\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_16\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_80\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_8\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_7\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_6\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_40\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_41\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_21\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_22\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_73\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_71\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_72\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_20\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_17\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_78\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_79\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_4\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_5\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_18\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_19\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_76\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_77\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_39\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_3\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_38\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_2\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_0\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_1\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_37\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_35\ : std_logic;
signal \switch_clk_1MHz_inst.current_stateZ0Z_1\ : std_logic;
signal \switch_clk_1MHz_inst_current_state_0\ : std_logic;
signal \switch_clk_1MHz_inst.bit_sequence_statZ0Z_36\ : std_logic;
signal \CLK_1_c_g\ : std_logic;
signal \switch_clk_1MHz_inst.N_377_g\ : std_logic;
signal \RST_N_c_i_g\ : std_logic;
signal \config_register_latched_dec_inst.STATCNF_0\ : std_logic;
signal \STATCNF_i_0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal xor_out_stat_wire : std_logic;
signal clk_output_wire : std_logic;
signal sel_output_wire : std_logic;
signal xor_out_dyn_wire : std_logic;
signal miso_input_wire : std_logic;
signal \RST_N_wire\ : std_logic;
signal mosi_output_wire : std_logic;
signal \CLK_wire\ : std_logic;

begin
    xor_out_stat <= xor_out_stat_wire;
    clk_output <= clk_output_wire;
    sel_output <= sel_output_wire;
    xor_out_dyn <= xor_out_dyn_wire;
    miso_input_wire <= miso_input;
    \RST_N_wire\ <= RST_N;
    mosi_output <= mosi_output_wire;
    \CLK_wire\ <= CLK;

    \xor_out_stat_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11095\,
            DIN => \N__11094\,
            DOUT => \N__11093\,
            PACKAGEPIN => xor_out_stat_wire
        );

    \xor_out_stat_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11095\,
            PADOUT => \N__11094\,
            PADIN => \N__11093\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9309\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11086\,
            DIN => \N__11085\,
            DOUT => \N__11084\,
            PACKAGEPIN => clk_output_wire
        );

    \clk_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11086\,
            PADOUT => \N__11085\,
            PADIN => \N__11084\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8439\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sel_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11077\,
            DIN => \N__11076\,
            DOUT => \N__11075\,
            PACKAGEPIN => sel_output_wire
        );

    \sel_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11077\,
            PADOUT => \N__11076\,
            PADIN => \N__11075\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8739\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \xor_out_dyn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11068\,
            DIN => \N__11067\,
            DOUT => \N__11066\,
            PACKAGEPIN => xor_out_dyn_wire
        );

    \xor_out_dyn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11068\,
            PADOUT => \N__11067\,
            PADIN => \N__11066\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5697\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \miso_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11059\,
            DIN => \N__11058\,
            DOUT => \N__11057\,
            PACKAGEPIN => miso_input_wire
        );

    \miso_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11059\,
            PADOUT => \N__11058\,
            PADIN => \N__11057\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => miso_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RST_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11050\,
            DIN => \N__11049\,
            DOUT => \N__11048\,
            PACKAGEPIN => \RST_N_wire\
        );

    \RST_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11050\,
            PADOUT => \N__11049\,
            PADIN => \N__11048\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RST_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \mosi_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11041\,
            DIN => \N__11040\,
            DOUT => \N__11039\,
            PACKAGEPIN => mosi_output_wire
        );

    \mosi_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11041\,
            PADOUT => \N__11040\,
            PADIN => \N__11039\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7197\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11032\,
            DIN => \N__11031\,
            DOUT => \N__11030\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11032\,
            PADOUT => \N__11031\,
            PADIN => \N__11030\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK_ibuf_gb_io_gb_input\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2561\ : InMux
    port map (
            O => \N__11013\,
            I => \N__11010\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__11010\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_38\
        );

    \I__2559\ : InMux
    port map (
            O => \N__11007\,
            I => \N__11004\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__11004\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_2\
        );

    \I__2557\ : InMux
    port map (
            O => \N__11001\,
            I => \N__10998\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__10998\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_0\
        );

    \I__2555\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10992\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__10992\,
            I => \N__10989\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__10989\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_1\
        );

    \I__2552\ : InMux
    port map (
            O => \N__10986\,
            I => \N__10983\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__10983\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_37\
        );

    \I__2550\ : InMux
    port map (
            O => \N__10980\,
            I => \N__10977\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__10977\,
            I => \N__10974\
        );

    \I__2548\ : Odrv12
    port map (
            O => \N__10974\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_35\
        );

    \I__2547\ : CascadeMux
    port map (
            O => \N__10971\,
            I => \N__10960\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__10970\,
            I => \N__10957\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__10969\,
            I => \N__10954\
        );

    \I__2544\ : CascadeMux
    port map (
            O => \N__10968\,
            I => \N__10951\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__10967\,
            I => \N__10931\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__10966\,
            I => \N__10928\
        );

    \I__2541\ : CascadeMux
    port map (
            O => \N__10965\,
            I => \N__10925\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__10964\,
            I => \N__10902\
        );

    \I__2539\ : CascadeMux
    port map (
            O => \N__10963\,
            I => \N__10899\
        );

    \I__2538\ : InMux
    port map (
            O => \N__10960\,
            I => \N__10861\
        );

    \I__2537\ : InMux
    port map (
            O => \N__10957\,
            I => \N__10861\
        );

    \I__2536\ : InMux
    port map (
            O => \N__10954\,
            I => \N__10861\
        );

    \I__2535\ : InMux
    port map (
            O => \N__10951\,
            I => \N__10861\
        );

    \I__2534\ : InMux
    port map (
            O => \N__10950\,
            I => \N__10861\
        );

    \I__2533\ : InMux
    port map (
            O => \N__10949\,
            I => \N__10861\
        );

    \I__2532\ : InMux
    port map (
            O => \N__10948\,
            I => \N__10861\
        );

    \I__2531\ : InMux
    port map (
            O => \N__10947\,
            I => \N__10852\
        );

    \I__2530\ : InMux
    port map (
            O => \N__10946\,
            I => \N__10852\
        );

    \I__2529\ : InMux
    port map (
            O => \N__10945\,
            I => \N__10852\
        );

    \I__2528\ : InMux
    port map (
            O => \N__10944\,
            I => \N__10852\
        );

    \I__2527\ : InMux
    port map (
            O => \N__10943\,
            I => \N__10847\
        );

    \I__2526\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10847\
        );

    \I__2525\ : InMux
    port map (
            O => \N__10941\,
            I => \N__10844\
        );

    \I__2524\ : InMux
    port map (
            O => \N__10940\,
            I => \N__10837\
        );

    \I__2523\ : InMux
    port map (
            O => \N__10939\,
            I => \N__10837\
        );

    \I__2522\ : InMux
    port map (
            O => \N__10938\,
            I => \N__10837\
        );

    \I__2521\ : InMux
    port map (
            O => \N__10937\,
            I => \N__10834\
        );

    \I__2520\ : InMux
    port map (
            O => \N__10936\,
            I => \N__10831\
        );

    \I__2519\ : InMux
    port map (
            O => \N__10935\,
            I => \N__10826\
        );

    \I__2518\ : InMux
    port map (
            O => \N__10934\,
            I => \N__10826\
        );

    \I__2517\ : InMux
    port map (
            O => \N__10931\,
            I => \N__10813\
        );

    \I__2516\ : InMux
    port map (
            O => \N__10928\,
            I => \N__10813\
        );

    \I__2515\ : InMux
    port map (
            O => \N__10925\,
            I => \N__10813\
        );

    \I__2514\ : InMux
    port map (
            O => \N__10924\,
            I => \N__10813\
        );

    \I__2513\ : InMux
    port map (
            O => \N__10923\,
            I => \N__10813\
        );

    \I__2512\ : InMux
    port map (
            O => \N__10922\,
            I => \N__10813\
        );

    \I__2511\ : InMux
    port map (
            O => \N__10921\,
            I => \N__10798\
        );

    \I__2510\ : InMux
    port map (
            O => \N__10920\,
            I => \N__10798\
        );

    \I__2509\ : InMux
    port map (
            O => \N__10919\,
            I => \N__10798\
        );

    \I__2508\ : InMux
    port map (
            O => \N__10918\,
            I => \N__10798\
        );

    \I__2507\ : InMux
    port map (
            O => \N__10917\,
            I => \N__10798\
        );

    \I__2506\ : InMux
    port map (
            O => \N__10916\,
            I => \N__10798\
        );

    \I__2505\ : InMux
    port map (
            O => \N__10915\,
            I => \N__10798\
        );

    \I__2504\ : InMux
    port map (
            O => \N__10914\,
            I => \N__10785\
        );

    \I__2503\ : InMux
    port map (
            O => \N__10913\,
            I => \N__10785\
        );

    \I__2502\ : InMux
    port map (
            O => \N__10912\,
            I => \N__10785\
        );

    \I__2501\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10785\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10910\,
            I => \N__10785\
        );

    \I__2499\ : InMux
    port map (
            O => \N__10909\,
            I => \N__10785\
        );

    \I__2498\ : InMux
    port map (
            O => \N__10908\,
            I => \N__10782\
        );

    \I__2497\ : InMux
    port map (
            O => \N__10907\,
            I => \N__10779\
        );

    \I__2496\ : InMux
    port map (
            O => \N__10906\,
            I => \N__10776\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10905\,
            I => \N__10773\
        );

    \I__2494\ : InMux
    port map (
            O => \N__10902\,
            I => \N__10742\
        );

    \I__2493\ : InMux
    port map (
            O => \N__10899\,
            I => \N__10742\
        );

    \I__2492\ : InMux
    port map (
            O => \N__10898\,
            I => \N__10742\
        );

    \I__2491\ : InMux
    port map (
            O => \N__10897\,
            I => \N__10742\
        );

    \I__2490\ : InMux
    port map (
            O => \N__10896\,
            I => \N__10742\
        );

    \I__2489\ : InMux
    port map (
            O => \N__10895\,
            I => \N__10742\
        );

    \I__2488\ : InMux
    port map (
            O => \N__10894\,
            I => \N__10742\
        );

    \I__2487\ : InMux
    port map (
            O => \N__10893\,
            I => \N__10737\
        );

    \I__2486\ : InMux
    port map (
            O => \N__10892\,
            I => \N__10737\
        );

    \I__2485\ : InMux
    port map (
            O => \N__10891\,
            I => \N__10734\
        );

    \I__2484\ : InMux
    port map (
            O => \N__10890\,
            I => \N__10731\
        );

    \I__2483\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10722\
        );

    \I__2482\ : InMux
    port map (
            O => \N__10888\,
            I => \N__10722\
        );

    \I__2481\ : InMux
    port map (
            O => \N__10887\,
            I => \N__10722\
        );

    \I__2480\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10722\
        );

    \I__2479\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10713\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10713\
        );

    \I__2477\ : InMux
    port map (
            O => \N__10883\,
            I => \N__10713\
        );

    \I__2476\ : InMux
    port map (
            O => \N__10882\,
            I => \N__10713\
        );

    \I__2475\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10700\
        );

    \I__2474\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10700\
        );

    \I__2473\ : InMux
    port map (
            O => \N__10879\,
            I => \N__10700\
        );

    \I__2472\ : InMux
    port map (
            O => \N__10878\,
            I => \N__10700\
        );

    \I__2471\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10700\
        );

    \I__2470\ : InMux
    port map (
            O => \N__10876\,
            I => \N__10700\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__10861\,
            I => \N__10693\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__10852\,
            I => \N__10693\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__10847\,
            I => \N__10693\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__10844\,
            I => \N__10688\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__10837\,
            I => \N__10688\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__10834\,
            I => \N__10683\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__10831\,
            I => \N__10683\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__10826\,
            I => \N__10675\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__10813\,
            I => \N__10668\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__10798\,
            I => \N__10668\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__10785\,
            I => \N__10668\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__10782\,
            I => \N__10659\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__10779\,
            I => \N__10659\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__10776\,
            I => \N__10659\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__10773\,
            I => \N__10659\
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__10772\,
            I => \N__10656\
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__10771\,
            I => \N__10642\
        );

    \I__2452\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10635\
        );

    \I__2451\ : InMux
    port map (
            O => \N__10769\,
            I => \N__10635\
        );

    \I__2450\ : InMux
    port map (
            O => \N__10768\,
            I => \N__10635\
        );

    \I__2449\ : InMux
    port map (
            O => \N__10767\,
            I => \N__10618\
        );

    \I__2448\ : InMux
    port map (
            O => \N__10766\,
            I => \N__10618\
        );

    \I__2447\ : InMux
    port map (
            O => \N__10765\,
            I => \N__10618\
        );

    \I__2446\ : InMux
    port map (
            O => \N__10764\,
            I => \N__10618\
        );

    \I__2445\ : InMux
    port map (
            O => \N__10763\,
            I => \N__10618\
        );

    \I__2444\ : InMux
    port map (
            O => \N__10762\,
            I => \N__10618\
        );

    \I__2443\ : InMux
    port map (
            O => \N__10761\,
            I => \N__10618\
        );

    \I__2442\ : InMux
    port map (
            O => \N__10760\,
            I => \N__10613\
        );

    \I__2441\ : InMux
    port map (
            O => \N__10759\,
            I => \N__10613\
        );

    \I__2440\ : InMux
    port map (
            O => \N__10758\,
            I => \N__10596\
        );

    \I__2439\ : InMux
    port map (
            O => \N__10757\,
            I => \N__10596\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__10742\,
            I => \N__10591\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__10737\,
            I => \N__10591\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__10734\,
            I => \N__10586\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__10731\,
            I => \N__10586\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__10722\,
            I => \N__10573\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__10713\,
            I => \N__10573\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__10700\,
            I => \N__10573\
        );

    \I__2431\ : Span4Mux_h
    port map (
            O => \N__10693\,
            I => \N__10573\
        );

    \I__2430\ : Span4Mux_v
    port map (
            O => \N__10688\,
            I => \N__10573\
        );

    \I__2429\ : Span4Mux_v
    port map (
            O => \N__10683\,
            I => \N__10573\
        );

    \I__2428\ : InMux
    port map (
            O => \N__10682\,
            I => \N__10566\
        );

    \I__2427\ : InMux
    port map (
            O => \N__10681\,
            I => \N__10566\
        );

    \I__2426\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10566\
        );

    \I__2425\ : InMux
    port map (
            O => \N__10679\,
            I => \N__10561\
        );

    \I__2424\ : InMux
    port map (
            O => \N__10678\,
            I => \N__10561\
        );

    \I__2423\ : Span4Mux_v
    port map (
            O => \N__10675\,
            I => \N__10554\
        );

    \I__2422\ : Span4Mux_v
    port map (
            O => \N__10668\,
            I => \N__10554\
        );

    \I__2421\ : Span4Mux_h
    port map (
            O => \N__10659\,
            I => \N__10554\
        );

    \I__2420\ : InMux
    port map (
            O => \N__10656\,
            I => \N__10549\
        );

    \I__2419\ : InMux
    port map (
            O => \N__10655\,
            I => \N__10549\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10654\,
            I => \N__10546\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10653\,
            I => \N__10537\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10652\,
            I => \N__10537\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10651\,
            I => \N__10537\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10650\,
            I => \N__10537\
        );

    \I__2413\ : InMux
    port map (
            O => \N__10649\,
            I => \N__10528\
        );

    \I__2412\ : InMux
    port map (
            O => \N__10648\,
            I => \N__10528\
        );

    \I__2411\ : InMux
    port map (
            O => \N__10647\,
            I => \N__10528\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10646\,
            I => \N__10528\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10645\,
            I => \N__10525\
        );

    \I__2408\ : InMux
    port map (
            O => \N__10642\,
            I => \N__10522\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__10635\,
            I => \N__10519\
        );

    \I__2406\ : InMux
    port map (
            O => \N__10634\,
            I => \N__10514\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10633\,
            I => \N__10514\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10618\,
            I => \N__10509\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__10613\,
            I => \N__10509\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__10612\,
            I => \N__10505\
        );

    \I__2401\ : InMux
    port map (
            O => \N__10611\,
            I => \N__10502\
        );

    \I__2400\ : InMux
    port map (
            O => \N__10610\,
            I => \N__10497\
        );

    \I__2399\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10497\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10608\,
            I => \N__10480\
        );

    \I__2397\ : InMux
    port map (
            O => \N__10607\,
            I => \N__10480\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10606\,
            I => \N__10480\
        );

    \I__2395\ : InMux
    port map (
            O => \N__10605\,
            I => \N__10480\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10604\,
            I => \N__10480\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10603\,
            I => \N__10480\
        );

    \I__2392\ : InMux
    port map (
            O => \N__10602\,
            I => \N__10480\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10480\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__10596\,
            I => \N__10477\
        );

    \I__2389\ : Span4Mux_v
    port map (
            O => \N__10591\,
            I => \N__10470\
        );

    \I__2388\ : Span4Mux_v
    port map (
            O => \N__10586\,
            I => \N__10470\
        );

    \I__2387\ : Span4Mux_h
    port map (
            O => \N__10573\,
            I => \N__10470\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__10566\,
            I => \N__10463\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__10561\,
            I => \N__10463\
        );

    \I__2384\ : Span4Mux_h
    port map (
            O => \N__10554\,
            I => \N__10463\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__10549\,
            I => \N__10458\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__10546\,
            I => \N__10458\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__10537\,
            I => \N__10443\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__10528\,
            I => \N__10443\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__10525\,
            I => \N__10443\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__10522\,
            I => \N__10443\
        );

    \I__2377\ : Span4Mux_v
    port map (
            O => \N__10519\,
            I => \N__10443\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__10514\,
            I => \N__10443\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__10509\,
            I => \N__10443\
        );

    \I__2374\ : InMux
    port map (
            O => \N__10508\,
            I => \N__10438\
        );

    \I__2373\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10438\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10502\,
            I => \switch_clk_1MHz_inst.current_stateZ0Z_1\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10497\,
            I => \switch_clk_1MHz_inst.current_stateZ0Z_1\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__10480\,
            I => \switch_clk_1MHz_inst.current_stateZ0Z_1\
        );

    \I__2369\ : Odrv12
    port map (
            O => \N__10477\,
            I => \switch_clk_1MHz_inst.current_stateZ0Z_1\
        );

    \I__2368\ : Odrv4
    port map (
            O => \N__10470\,
            I => \switch_clk_1MHz_inst.current_stateZ0Z_1\
        );

    \I__2367\ : Odrv4
    port map (
            O => \N__10463\,
            I => \switch_clk_1MHz_inst.current_stateZ0Z_1\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__10458\,
            I => \switch_clk_1MHz_inst.current_stateZ0Z_1\
        );

    \I__2365\ : Odrv4
    port map (
            O => \N__10443\,
            I => \switch_clk_1MHz_inst.current_stateZ0Z_1\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__10438\,
            I => \switch_clk_1MHz_inst.current_stateZ0Z_1\
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__10419\,
            I => \N__10405\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__10418\,
            I => \N__10400\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__10417\,
            I => \N__10397\
        );

    \I__2360\ : CascadeMux
    port map (
            O => \N__10416\,
            I => \N__10394\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__10415\,
            I => \N__10391\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10414\,
            I => \N__10369\
        );

    \I__2357\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10364\
        );

    \I__2356\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10364\
        );

    \I__2355\ : CascadeMux
    port map (
            O => \N__10411\,
            I => \N__10360\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__10410\,
            I => \N__10357\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__10409\,
            I => \N__10354\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__10408\,
            I => \N__10344\
        );

    \I__2351\ : InMux
    port map (
            O => \N__10405\,
            I => \N__10336\
        );

    \I__2350\ : InMux
    port map (
            O => \N__10404\,
            I => \N__10336\
        );

    \I__2349\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10336\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10321\
        );

    \I__2347\ : InMux
    port map (
            O => \N__10397\,
            I => \N__10321\
        );

    \I__2346\ : InMux
    port map (
            O => \N__10394\,
            I => \N__10321\
        );

    \I__2345\ : InMux
    port map (
            O => \N__10391\,
            I => \N__10321\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10390\,
            I => \N__10321\
        );

    \I__2343\ : InMux
    port map (
            O => \N__10389\,
            I => \N__10321\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10388\,
            I => \N__10321\
        );

    \I__2341\ : InMux
    port map (
            O => \N__10387\,
            I => \N__10313\
        );

    \I__2340\ : InMux
    port map (
            O => \N__10386\,
            I => \N__10313\
        );

    \I__2339\ : InMux
    port map (
            O => \N__10385\,
            I => \N__10310\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__10384\,
            I => \N__10305\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__10383\,
            I => \N__10302\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__10382\,
            I => \N__10299\
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__10381\,
            I => \N__10296\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__10380\,
            I => \N__10291\
        );

    \I__2333\ : InMux
    port map (
            O => \N__10379\,
            I => \N__10286\
        );

    \I__2332\ : InMux
    port map (
            O => \N__10378\,
            I => \N__10273\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10377\,
            I => \N__10273\
        );

    \I__2330\ : InMux
    port map (
            O => \N__10376\,
            I => \N__10273\
        );

    \I__2329\ : InMux
    port map (
            O => \N__10375\,
            I => \N__10273\
        );

    \I__2328\ : InMux
    port map (
            O => \N__10374\,
            I => \N__10273\
        );

    \I__2327\ : InMux
    port map (
            O => \N__10373\,
            I => \N__10273\
        );

    \I__2326\ : InMux
    port map (
            O => \N__10372\,
            I => \N__10270\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__10369\,
            I => \N__10265\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__10364\,
            I => \N__10265\
        );

    \I__2323\ : InMux
    port map (
            O => \N__10363\,
            I => \N__10255\
        );

    \I__2322\ : InMux
    port map (
            O => \N__10360\,
            I => \N__10242\
        );

    \I__2321\ : InMux
    port map (
            O => \N__10357\,
            I => \N__10242\
        );

    \I__2320\ : InMux
    port map (
            O => \N__10354\,
            I => \N__10242\
        );

    \I__2319\ : InMux
    port map (
            O => \N__10353\,
            I => \N__10242\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10352\,
            I => \N__10242\
        );

    \I__2317\ : InMux
    port map (
            O => \N__10351\,
            I => \N__10242\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__10350\,
            I => \N__10239\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__10349\,
            I => \N__10236\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__10348\,
            I => \N__10233\
        );

    \I__2313\ : CascadeMux
    port map (
            O => \N__10347\,
            I => \N__10230\
        );

    \I__2312\ : InMux
    port map (
            O => \N__10344\,
            I => \N__10184\
        );

    \I__2311\ : InMux
    port map (
            O => \N__10343\,
            I => \N__10184\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__10336\,
            I => \N__10179\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__10321\,
            I => \N__10179\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10320\,
            I => \N__10174\
        );

    \I__2307\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10174\
        );

    \I__2306\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10171\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__10313\,
            I => \N__10166\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__10310\,
            I => \N__10166\
        );

    \I__2303\ : InMux
    port map (
            O => \N__10309\,
            I => \N__10151\
        );

    \I__2302\ : InMux
    port map (
            O => \N__10308\,
            I => \N__10151\
        );

    \I__2301\ : InMux
    port map (
            O => \N__10305\,
            I => \N__10151\
        );

    \I__2300\ : InMux
    port map (
            O => \N__10302\,
            I => \N__10151\
        );

    \I__2299\ : InMux
    port map (
            O => \N__10299\,
            I => \N__10151\
        );

    \I__2298\ : InMux
    port map (
            O => \N__10296\,
            I => \N__10151\
        );

    \I__2297\ : InMux
    port map (
            O => \N__10295\,
            I => \N__10151\
        );

    \I__2296\ : InMux
    port map (
            O => \N__10294\,
            I => \N__10148\
        );

    \I__2295\ : InMux
    port map (
            O => \N__10291\,
            I => \N__10141\
        );

    \I__2294\ : InMux
    port map (
            O => \N__10290\,
            I => \N__10141\
        );

    \I__2293\ : InMux
    port map (
            O => \N__10289\,
            I => \N__10141\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__10286\,
            I => \N__10136\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__10273\,
            I => \N__10136\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__10270\,
            I => \N__10131\
        );

    \I__2289\ : Span4Mux_v
    port map (
            O => \N__10265\,
            I => \N__10131\
        );

    \I__2288\ : InMux
    port map (
            O => \N__10264\,
            I => \N__10128\
        );

    \I__2287\ : InMux
    port map (
            O => \N__10263\,
            I => \N__10121\
        );

    \I__2286\ : InMux
    port map (
            O => \N__10262\,
            I => \N__10121\
        );

    \I__2285\ : InMux
    port map (
            O => \N__10261\,
            I => \N__10121\
        );

    \I__2284\ : InMux
    port map (
            O => \N__10260\,
            I => \N__10114\
        );

    \I__2283\ : InMux
    port map (
            O => \N__10259\,
            I => \N__10114\
        );

    \I__2282\ : InMux
    port map (
            O => \N__10258\,
            I => \N__10114\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__10255\,
            I => \N__10109\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__10242\,
            I => \N__10109\
        );

    \I__2279\ : InMux
    port map (
            O => \N__10239\,
            I => \N__10082\
        );

    \I__2278\ : InMux
    port map (
            O => \N__10236\,
            I => \N__10082\
        );

    \I__2277\ : InMux
    port map (
            O => \N__10233\,
            I => \N__10082\
        );

    \I__2276\ : InMux
    port map (
            O => \N__10230\,
            I => \N__10082\
        );

    \I__2275\ : InMux
    port map (
            O => \N__10229\,
            I => \N__10082\
        );

    \I__2274\ : InMux
    port map (
            O => \N__10228\,
            I => \N__10082\
        );

    \I__2273\ : InMux
    port map (
            O => \N__10227\,
            I => \N__10082\
        );

    \I__2272\ : InMux
    port map (
            O => \N__10226\,
            I => \N__10077\
        );

    \I__2271\ : InMux
    port map (
            O => \N__10225\,
            I => \N__10077\
        );

    \I__2270\ : InMux
    port map (
            O => \N__10224\,
            I => \N__10072\
        );

    \I__2269\ : InMux
    port map (
            O => \N__10223\,
            I => \N__10072\
        );

    \I__2268\ : InMux
    port map (
            O => \N__10222\,
            I => \N__10063\
        );

    \I__2267\ : InMux
    port map (
            O => \N__10221\,
            I => \N__10063\
        );

    \I__2266\ : InMux
    port map (
            O => \N__10220\,
            I => \N__10063\
        );

    \I__2265\ : InMux
    port map (
            O => \N__10219\,
            I => \N__10063\
        );

    \I__2264\ : InMux
    port map (
            O => \N__10218\,
            I => \N__10060\
        );

    \I__2263\ : InMux
    port map (
            O => \N__10217\,
            I => \N__10055\
        );

    \I__2262\ : InMux
    port map (
            O => \N__10216\,
            I => \N__10055\
        );

    \I__2261\ : InMux
    port map (
            O => \N__10215\,
            I => \N__10050\
        );

    \I__2260\ : InMux
    port map (
            O => \N__10214\,
            I => \N__10050\
        );

    \I__2259\ : InMux
    port map (
            O => \N__10213\,
            I => \N__10035\
        );

    \I__2258\ : InMux
    port map (
            O => \N__10212\,
            I => \N__10035\
        );

    \I__2257\ : InMux
    port map (
            O => \N__10211\,
            I => \N__10035\
        );

    \I__2256\ : InMux
    port map (
            O => \N__10210\,
            I => \N__10035\
        );

    \I__2255\ : InMux
    port map (
            O => \N__10209\,
            I => \N__10035\
        );

    \I__2254\ : InMux
    port map (
            O => \N__10208\,
            I => \N__10035\
        );

    \I__2253\ : InMux
    port map (
            O => \N__10207\,
            I => \N__10035\
        );

    \I__2252\ : InMux
    port map (
            O => \N__10206\,
            I => \N__10018\
        );

    \I__2251\ : InMux
    port map (
            O => \N__10205\,
            I => \N__10018\
        );

    \I__2250\ : InMux
    port map (
            O => \N__10204\,
            I => \N__10018\
        );

    \I__2249\ : InMux
    port map (
            O => \N__10203\,
            I => \N__10018\
        );

    \I__2248\ : InMux
    port map (
            O => \N__10202\,
            I => \N__10018\
        );

    \I__2247\ : InMux
    port map (
            O => \N__10201\,
            I => \N__10018\
        );

    \I__2246\ : InMux
    port map (
            O => \N__10200\,
            I => \N__10018\
        );

    \I__2245\ : InMux
    port map (
            O => \N__10199\,
            I => \N__10018\
        );

    \I__2244\ : InMux
    port map (
            O => \N__10198\,
            I => \N__10001\
        );

    \I__2243\ : InMux
    port map (
            O => \N__10197\,
            I => \N__10001\
        );

    \I__2242\ : InMux
    port map (
            O => \N__10196\,
            I => \N__10001\
        );

    \I__2241\ : InMux
    port map (
            O => \N__10195\,
            I => \N__10001\
        );

    \I__2240\ : InMux
    port map (
            O => \N__10194\,
            I => \N__10001\
        );

    \I__2239\ : InMux
    port map (
            O => \N__10193\,
            I => \N__10001\
        );

    \I__2238\ : InMux
    port map (
            O => \N__10192\,
            I => \N__10001\
        );

    \I__2237\ : InMux
    port map (
            O => \N__10191\,
            I => \N__10001\
        );

    \I__2236\ : InMux
    port map (
            O => \N__10190\,
            I => \N__9993\
        );

    \I__2235\ : InMux
    port map (
            O => \N__10189\,
            I => \N__9993\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__10184\,
            I => \N__9990\
        );

    \I__2233\ : Span4Mux_h
    port map (
            O => \N__10179\,
            I => \N__9987\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__10174\,
            I => \N__9980\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__10171\,
            I => \N__9980\
        );

    \I__2230\ : Span4Mux_h
    port map (
            O => \N__10166\,
            I => \N__9980\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__10151\,
            I => \N__9976\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__10148\,
            I => \N__9969\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__10141\,
            I => \N__9969\
        );

    \I__2226\ : Span4Mux_h
    port map (
            O => \N__10136\,
            I => \N__9969\
        );

    \I__2225\ : Span4Mux_h
    port map (
            O => \N__10131\,
            I => \N__9964\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__10128\,
            I => \N__9964\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__10121\,
            I => \N__9957\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__10114\,
            I => \N__9957\
        );

    \I__2221\ : Span4Mux_h
    port map (
            O => \N__10109\,
            I => \N__9957\
        );

    \I__2220\ : InMux
    port map (
            O => \N__10108\,
            I => \N__9948\
        );

    \I__2219\ : InMux
    port map (
            O => \N__10107\,
            I => \N__9948\
        );

    \I__2218\ : InMux
    port map (
            O => \N__10106\,
            I => \N__9948\
        );

    \I__2217\ : InMux
    port map (
            O => \N__10105\,
            I => \N__9948\
        );

    \I__2216\ : InMux
    port map (
            O => \N__10104\,
            I => \N__9935\
        );

    \I__2215\ : InMux
    port map (
            O => \N__10103\,
            I => \N__9935\
        );

    \I__2214\ : InMux
    port map (
            O => \N__10102\,
            I => \N__9935\
        );

    \I__2213\ : InMux
    port map (
            O => \N__10101\,
            I => \N__9935\
        );

    \I__2212\ : InMux
    port map (
            O => \N__10100\,
            I => \N__9926\
        );

    \I__2211\ : InMux
    port map (
            O => \N__10099\,
            I => \N__9926\
        );

    \I__2210\ : InMux
    port map (
            O => \N__10098\,
            I => \N__9926\
        );

    \I__2209\ : InMux
    port map (
            O => \N__10097\,
            I => \N__9926\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__10082\,
            I => \N__9923\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__10077\,
            I => \N__9904\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__10072\,
            I => \N__9904\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__10063\,
            I => \N__9904\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__10060\,
            I => \N__9904\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__10055\,
            I => \N__9904\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__10050\,
            I => \N__9904\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__10035\,
            I => \N__9904\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__10018\,
            I => \N__9904\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__10001\,
            I => \N__9904\
        );

    \I__2198\ : InMux
    port map (
            O => \N__10000\,
            I => \N__9899\
        );

    \I__2197\ : InMux
    port map (
            O => \N__9999\,
            I => \N__9899\
        );

    \I__2196\ : InMux
    port map (
            O => \N__9998\,
            I => \N__9896\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__9993\,
            I => \N__9887\
        );

    \I__2194\ : Span4Mux_s3_h
    port map (
            O => \N__9990\,
            I => \N__9887\
        );

    \I__2193\ : Span4Mux_h
    port map (
            O => \N__9987\,
            I => \N__9887\
        );

    \I__2192\ : Span4Mux_h
    port map (
            O => \N__9980\,
            I => \N__9887\
        );

    \I__2191\ : InMux
    port map (
            O => \N__9979\,
            I => \N__9884\
        );

    \I__2190\ : Span4Mux_s3_h
    port map (
            O => \N__9976\,
            I => \N__9877\
        );

    \I__2189\ : Span4Mux_h
    port map (
            O => \N__9969\,
            I => \N__9877\
        );

    \I__2188\ : Span4Mux_h
    port map (
            O => \N__9964\,
            I => \N__9877\
        );

    \I__2187\ : Span4Mux_h
    port map (
            O => \N__9957\,
            I => \N__9872\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9948\,
            I => \N__9872\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9947\,
            I => \N__9863\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9863\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9863\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9944\,
            I => \N__9863\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9935\,
            I => \switch_clk_1MHz_inst_current_state_0\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__9926\,
            I => \switch_clk_1MHz_inst_current_state_0\
        );

    \I__2179\ : Odrv4
    port map (
            O => \N__9923\,
            I => \switch_clk_1MHz_inst_current_state_0\
        );

    \I__2178\ : Odrv12
    port map (
            O => \N__9904\,
            I => \switch_clk_1MHz_inst_current_state_0\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__9899\,
            I => \switch_clk_1MHz_inst_current_state_0\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9896\,
            I => \switch_clk_1MHz_inst_current_state_0\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__9887\,
            I => \switch_clk_1MHz_inst_current_state_0\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__9884\,
            I => \switch_clk_1MHz_inst_current_state_0\
        );

    \I__2173\ : Odrv4
    port map (
            O => \N__9877\,
            I => \switch_clk_1MHz_inst_current_state_0\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__9872\,
            I => \switch_clk_1MHz_inst_current_state_0\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__9863\,
            I => \switch_clk_1MHz_inst_current_state_0\
        );

    \I__2170\ : InMux
    port map (
            O => \N__9840\,
            I => \N__9837\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__9837\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_36\
        );

    \I__2168\ : ClkMux
    port map (
            O => \N__9834\,
            I => \N__9624\
        );

    \I__2167\ : ClkMux
    port map (
            O => \N__9833\,
            I => \N__9624\
        );

    \I__2166\ : ClkMux
    port map (
            O => \N__9832\,
            I => \N__9624\
        );

    \I__2165\ : ClkMux
    port map (
            O => \N__9831\,
            I => \N__9624\
        );

    \I__2164\ : ClkMux
    port map (
            O => \N__9830\,
            I => \N__9624\
        );

    \I__2163\ : ClkMux
    port map (
            O => \N__9829\,
            I => \N__9624\
        );

    \I__2162\ : ClkMux
    port map (
            O => \N__9828\,
            I => \N__9624\
        );

    \I__2161\ : ClkMux
    port map (
            O => \N__9827\,
            I => \N__9624\
        );

    \I__2160\ : ClkMux
    port map (
            O => \N__9826\,
            I => \N__9624\
        );

    \I__2159\ : ClkMux
    port map (
            O => \N__9825\,
            I => \N__9624\
        );

    \I__2158\ : ClkMux
    port map (
            O => \N__9824\,
            I => \N__9624\
        );

    \I__2157\ : ClkMux
    port map (
            O => \N__9823\,
            I => \N__9624\
        );

    \I__2156\ : ClkMux
    port map (
            O => \N__9822\,
            I => \N__9624\
        );

    \I__2155\ : ClkMux
    port map (
            O => \N__9821\,
            I => \N__9624\
        );

    \I__2154\ : ClkMux
    port map (
            O => \N__9820\,
            I => \N__9624\
        );

    \I__2153\ : ClkMux
    port map (
            O => \N__9819\,
            I => \N__9624\
        );

    \I__2152\ : ClkMux
    port map (
            O => \N__9818\,
            I => \N__9624\
        );

    \I__2151\ : ClkMux
    port map (
            O => \N__9817\,
            I => \N__9624\
        );

    \I__2150\ : ClkMux
    port map (
            O => \N__9816\,
            I => \N__9624\
        );

    \I__2149\ : ClkMux
    port map (
            O => \N__9815\,
            I => \N__9624\
        );

    \I__2148\ : ClkMux
    port map (
            O => \N__9814\,
            I => \N__9624\
        );

    \I__2147\ : ClkMux
    port map (
            O => \N__9813\,
            I => \N__9624\
        );

    \I__2146\ : ClkMux
    port map (
            O => \N__9812\,
            I => \N__9624\
        );

    \I__2145\ : ClkMux
    port map (
            O => \N__9811\,
            I => \N__9624\
        );

    \I__2144\ : ClkMux
    port map (
            O => \N__9810\,
            I => \N__9624\
        );

    \I__2143\ : ClkMux
    port map (
            O => \N__9809\,
            I => \N__9624\
        );

    \I__2142\ : ClkMux
    port map (
            O => \N__9808\,
            I => \N__9624\
        );

    \I__2141\ : ClkMux
    port map (
            O => \N__9807\,
            I => \N__9624\
        );

    \I__2140\ : ClkMux
    port map (
            O => \N__9806\,
            I => \N__9624\
        );

    \I__2139\ : ClkMux
    port map (
            O => \N__9805\,
            I => \N__9624\
        );

    \I__2138\ : ClkMux
    port map (
            O => \N__9804\,
            I => \N__9624\
        );

    \I__2137\ : ClkMux
    port map (
            O => \N__9803\,
            I => \N__9624\
        );

    \I__2136\ : ClkMux
    port map (
            O => \N__9802\,
            I => \N__9624\
        );

    \I__2135\ : ClkMux
    port map (
            O => \N__9801\,
            I => \N__9624\
        );

    \I__2134\ : ClkMux
    port map (
            O => \N__9800\,
            I => \N__9624\
        );

    \I__2133\ : ClkMux
    port map (
            O => \N__9799\,
            I => \N__9624\
        );

    \I__2132\ : ClkMux
    port map (
            O => \N__9798\,
            I => \N__9624\
        );

    \I__2131\ : ClkMux
    port map (
            O => \N__9797\,
            I => \N__9624\
        );

    \I__2130\ : ClkMux
    port map (
            O => \N__9796\,
            I => \N__9624\
        );

    \I__2129\ : ClkMux
    port map (
            O => \N__9795\,
            I => \N__9624\
        );

    \I__2128\ : ClkMux
    port map (
            O => \N__9794\,
            I => \N__9624\
        );

    \I__2127\ : ClkMux
    port map (
            O => \N__9793\,
            I => \N__9624\
        );

    \I__2126\ : ClkMux
    port map (
            O => \N__9792\,
            I => \N__9624\
        );

    \I__2125\ : ClkMux
    port map (
            O => \N__9791\,
            I => \N__9624\
        );

    \I__2124\ : ClkMux
    port map (
            O => \N__9790\,
            I => \N__9624\
        );

    \I__2123\ : ClkMux
    port map (
            O => \N__9789\,
            I => \N__9624\
        );

    \I__2122\ : ClkMux
    port map (
            O => \N__9788\,
            I => \N__9624\
        );

    \I__2121\ : ClkMux
    port map (
            O => \N__9787\,
            I => \N__9624\
        );

    \I__2120\ : ClkMux
    port map (
            O => \N__9786\,
            I => \N__9624\
        );

    \I__2119\ : ClkMux
    port map (
            O => \N__9785\,
            I => \N__9624\
        );

    \I__2118\ : ClkMux
    port map (
            O => \N__9784\,
            I => \N__9624\
        );

    \I__2117\ : ClkMux
    port map (
            O => \N__9783\,
            I => \N__9624\
        );

    \I__2116\ : ClkMux
    port map (
            O => \N__9782\,
            I => \N__9624\
        );

    \I__2115\ : ClkMux
    port map (
            O => \N__9781\,
            I => \N__9624\
        );

    \I__2114\ : ClkMux
    port map (
            O => \N__9780\,
            I => \N__9624\
        );

    \I__2113\ : ClkMux
    port map (
            O => \N__9779\,
            I => \N__9624\
        );

    \I__2112\ : ClkMux
    port map (
            O => \N__9778\,
            I => \N__9624\
        );

    \I__2111\ : ClkMux
    port map (
            O => \N__9777\,
            I => \N__9624\
        );

    \I__2110\ : ClkMux
    port map (
            O => \N__9776\,
            I => \N__9624\
        );

    \I__2109\ : ClkMux
    port map (
            O => \N__9775\,
            I => \N__9624\
        );

    \I__2108\ : ClkMux
    port map (
            O => \N__9774\,
            I => \N__9624\
        );

    \I__2107\ : ClkMux
    port map (
            O => \N__9773\,
            I => \N__9624\
        );

    \I__2106\ : ClkMux
    port map (
            O => \N__9772\,
            I => \N__9624\
        );

    \I__2105\ : ClkMux
    port map (
            O => \N__9771\,
            I => \N__9624\
        );

    \I__2104\ : ClkMux
    port map (
            O => \N__9770\,
            I => \N__9624\
        );

    \I__2103\ : ClkMux
    port map (
            O => \N__9769\,
            I => \N__9624\
        );

    \I__2102\ : ClkMux
    port map (
            O => \N__9768\,
            I => \N__9624\
        );

    \I__2101\ : ClkMux
    port map (
            O => \N__9767\,
            I => \N__9624\
        );

    \I__2100\ : ClkMux
    port map (
            O => \N__9766\,
            I => \N__9624\
        );

    \I__2099\ : ClkMux
    port map (
            O => \N__9765\,
            I => \N__9624\
        );

    \I__2098\ : GlobalMux
    port map (
            O => \N__9624\,
            I => \N__9621\
        );

    \I__2097\ : gio2CtrlBuf
    port map (
            O => \N__9621\,
            I => \CLK_1_c_g\
        );

    \I__2096\ : CEMux
    port map (
            O => \N__9618\,
            I => \N__9546\
        );

    \I__2095\ : CEMux
    port map (
            O => \N__9617\,
            I => \N__9546\
        );

    \I__2094\ : CEMux
    port map (
            O => \N__9616\,
            I => \N__9546\
        );

    \I__2093\ : CEMux
    port map (
            O => \N__9615\,
            I => \N__9546\
        );

    \I__2092\ : CEMux
    port map (
            O => \N__9614\,
            I => \N__9546\
        );

    \I__2091\ : CEMux
    port map (
            O => \N__9613\,
            I => \N__9546\
        );

    \I__2090\ : CEMux
    port map (
            O => \N__9612\,
            I => \N__9546\
        );

    \I__2089\ : CEMux
    port map (
            O => \N__9611\,
            I => \N__9546\
        );

    \I__2088\ : CEMux
    port map (
            O => \N__9610\,
            I => \N__9546\
        );

    \I__2087\ : CEMux
    port map (
            O => \N__9609\,
            I => \N__9546\
        );

    \I__2086\ : CEMux
    port map (
            O => \N__9608\,
            I => \N__9546\
        );

    \I__2085\ : CEMux
    port map (
            O => \N__9607\,
            I => \N__9546\
        );

    \I__2084\ : CEMux
    port map (
            O => \N__9606\,
            I => \N__9546\
        );

    \I__2083\ : CEMux
    port map (
            O => \N__9605\,
            I => \N__9546\
        );

    \I__2082\ : CEMux
    port map (
            O => \N__9604\,
            I => \N__9546\
        );

    \I__2081\ : CEMux
    port map (
            O => \N__9603\,
            I => \N__9546\
        );

    \I__2080\ : CEMux
    port map (
            O => \N__9602\,
            I => \N__9546\
        );

    \I__2079\ : CEMux
    port map (
            O => \N__9601\,
            I => \N__9546\
        );

    \I__2078\ : CEMux
    port map (
            O => \N__9600\,
            I => \N__9546\
        );

    \I__2077\ : CEMux
    port map (
            O => \N__9599\,
            I => \N__9546\
        );

    \I__2076\ : CEMux
    port map (
            O => \N__9598\,
            I => \N__9546\
        );

    \I__2075\ : CEMux
    port map (
            O => \N__9597\,
            I => \N__9546\
        );

    \I__2074\ : CEMux
    port map (
            O => \N__9596\,
            I => \N__9546\
        );

    \I__2073\ : CEMux
    port map (
            O => \N__9595\,
            I => \N__9546\
        );

    \I__2072\ : GlobalMux
    port map (
            O => \N__9546\,
            I => \N__9543\
        );

    \I__2071\ : gio2CtrlBuf
    port map (
            O => \N__9543\,
            I => \switch_clk_1MHz_inst.N_377_g\
        );

    \I__2070\ : SRMux
    port map (
            O => \N__9540\,
            I => \N__9330\
        );

    \I__2069\ : SRMux
    port map (
            O => \N__9539\,
            I => \N__9330\
        );

    \I__2068\ : SRMux
    port map (
            O => \N__9538\,
            I => \N__9330\
        );

    \I__2067\ : SRMux
    port map (
            O => \N__9537\,
            I => \N__9330\
        );

    \I__2066\ : SRMux
    port map (
            O => \N__9536\,
            I => \N__9330\
        );

    \I__2065\ : SRMux
    port map (
            O => \N__9535\,
            I => \N__9330\
        );

    \I__2064\ : SRMux
    port map (
            O => \N__9534\,
            I => \N__9330\
        );

    \I__2063\ : SRMux
    port map (
            O => \N__9533\,
            I => \N__9330\
        );

    \I__2062\ : SRMux
    port map (
            O => \N__9532\,
            I => \N__9330\
        );

    \I__2061\ : SRMux
    port map (
            O => \N__9531\,
            I => \N__9330\
        );

    \I__2060\ : SRMux
    port map (
            O => \N__9530\,
            I => \N__9330\
        );

    \I__2059\ : SRMux
    port map (
            O => \N__9529\,
            I => \N__9330\
        );

    \I__2058\ : SRMux
    port map (
            O => \N__9528\,
            I => \N__9330\
        );

    \I__2057\ : SRMux
    port map (
            O => \N__9527\,
            I => \N__9330\
        );

    \I__2056\ : SRMux
    port map (
            O => \N__9526\,
            I => \N__9330\
        );

    \I__2055\ : SRMux
    port map (
            O => \N__9525\,
            I => \N__9330\
        );

    \I__2054\ : SRMux
    port map (
            O => \N__9524\,
            I => \N__9330\
        );

    \I__2053\ : SRMux
    port map (
            O => \N__9523\,
            I => \N__9330\
        );

    \I__2052\ : SRMux
    port map (
            O => \N__9522\,
            I => \N__9330\
        );

    \I__2051\ : SRMux
    port map (
            O => \N__9521\,
            I => \N__9330\
        );

    \I__2050\ : SRMux
    port map (
            O => \N__9520\,
            I => \N__9330\
        );

    \I__2049\ : SRMux
    port map (
            O => \N__9519\,
            I => \N__9330\
        );

    \I__2048\ : SRMux
    port map (
            O => \N__9518\,
            I => \N__9330\
        );

    \I__2047\ : SRMux
    port map (
            O => \N__9517\,
            I => \N__9330\
        );

    \I__2046\ : SRMux
    port map (
            O => \N__9516\,
            I => \N__9330\
        );

    \I__2045\ : SRMux
    port map (
            O => \N__9515\,
            I => \N__9330\
        );

    \I__2044\ : SRMux
    port map (
            O => \N__9514\,
            I => \N__9330\
        );

    \I__2043\ : SRMux
    port map (
            O => \N__9513\,
            I => \N__9330\
        );

    \I__2042\ : SRMux
    port map (
            O => \N__9512\,
            I => \N__9330\
        );

    \I__2041\ : SRMux
    port map (
            O => \N__9511\,
            I => \N__9330\
        );

    \I__2040\ : SRMux
    port map (
            O => \N__9510\,
            I => \N__9330\
        );

    \I__2039\ : SRMux
    port map (
            O => \N__9509\,
            I => \N__9330\
        );

    \I__2038\ : SRMux
    port map (
            O => \N__9508\,
            I => \N__9330\
        );

    \I__2037\ : SRMux
    port map (
            O => \N__9507\,
            I => \N__9330\
        );

    \I__2036\ : SRMux
    port map (
            O => \N__9506\,
            I => \N__9330\
        );

    \I__2035\ : SRMux
    port map (
            O => \N__9505\,
            I => \N__9330\
        );

    \I__2034\ : SRMux
    port map (
            O => \N__9504\,
            I => \N__9330\
        );

    \I__2033\ : SRMux
    port map (
            O => \N__9503\,
            I => \N__9330\
        );

    \I__2032\ : SRMux
    port map (
            O => \N__9502\,
            I => \N__9330\
        );

    \I__2031\ : SRMux
    port map (
            O => \N__9501\,
            I => \N__9330\
        );

    \I__2030\ : SRMux
    port map (
            O => \N__9500\,
            I => \N__9330\
        );

    \I__2029\ : SRMux
    port map (
            O => \N__9499\,
            I => \N__9330\
        );

    \I__2028\ : SRMux
    port map (
            O => \N__9498\,
            I => \N__9330\
        );

    \I__2027\ : SRMux
    port map (
            O => \N__9497\,
            I => \N__9330\
        );

    \I__2026\ : SRMux
    port map (
            O => \N__9496\,
            I => \N__9330\
        );

    \I__2025\ : SRMux
    port map (
            O => \N__9495\,
            I => \N__9330\
        );

    \I__2024\ : SRMux
    port map (
            O => \N__9494\,
            I => \N__9330\
        );

    \I__2023\ : SRMux
    port map (
            O => \N__9493\,
            I => \N__9330\
        );

    \I__2022\ : SRMux
    port map (
            O => \N__9492\,
            I => \N__9330\
        );

    \I__2021\ : SRMux
    port map (
            O => \N__9491\,
            I => \N__9330\
        );

    \I__2020\ : SRMux
    port map (
            O => \N__9490\,
            I => \N__9330\
        );

    \I__2019\ : SRMux
    port map (
            O => \N__9489\,
            I => \N__9330\
        );

    \I__2018\ : SRMux
    port map (
            O => \N__9488\,
            I => \N__9330\
        );

    \I__2017\ : SRMux
    port map (
            O => \N__9487\,
            I => \N__9330\
        );

    \I__2016\ : SRMux
    port map (
            O => \N__9486\,
            I => \N__9330\
        );

    \I__2015\ : SRMux
    port map (
            O => \N__9485\,
            I => \N__9330\
        );

    \I__2014\ : SRMux
    port map (
            O => \N__9484\,
            I => \N__9330\
        );

    \I__2013\ : SRMux
    port map (
            O => \N__9483\,
            I => \N__9330\
        );

    \I__2012\ : SRMux
    port map (
            O => \N__9482\,
            I => \N__9330\
        );

    \I__2011\ : SRMux
    port map (
            O => \N__9481\,
            I => \N__9330\
        );

    \I__2010\ : SRMux
    port map (
            O => \N__9480\,
            I => \N__9330\
        );

    \I__2009\ : SRMux
    port map (
            O => \N__9479\,
            I => \N__9330\
        );

    \I__2008\ : SRMux
    port map (
            O => \N__9478\,
            I => \N__9330\
        );

    \I__2007\ : SRMux
    port map (
            O => \N__9477\,
            I => \N__9330\
        );

    \I__2006\ : SRMux
    port map (
            O => \N__9476\,
            I => \N__9330\
        );

    \I__2005\ : SRMux
    port map (
            O => \N__9475\,
            I => \N__9330\
        );

    \I__2004\ : SRMux
    port map (
            O => \N__9474\,
            I => \N__9330\
        );

    \I__2003\ : SRMux
    port map (
            O => \N__9473\,
            I => \N__9330\
        );

    \I__2002\ : SRMux
    port map (
            O => \N__9472\,
            I => \N__9330\
        );

    \I__2001\ : SRMux
    port map (
            O => \N__9471\,
            I => \N__9330\
        );

    \I__2000\ : GlobalMux
    port map (
            O => \N__9330\,
            I => \N__9327\
        );

    \I__1999\ : gio2CtrlBuf
    port map (
            O => \N__9327\,
            I => \RST_N_c_i_g\
        );

    \I__1998\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9321\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__9321\,
            I => \N__9318\
        );

    \I__1996\ : Span12Mux_s2_h
    port map (
            O => \N__9318\,
            I => \N__9315\
        );

    \I__1995\ : Span12Mux_h
    port map (
            O => \N__9315\,
            I => \N__9312\
        );

    \I__1994\ : Odrv12
    port map (
            O => \N__9312\,
            I => \config_register_latched_dec_inst.STATCNF_0\
        );

    \I__1993\ : IoInMux
    port map (
            O => \N__9309\,
            I => \N__9306\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__9306\,
            I => \STATCNF_i_0\
        );

    \I__1991\ : InMux
    port map (
            O => \N__9303\,
            I => \N__9300\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__9300\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_17\
        );

    \I__1989\ : InMux
    port map (
            O => \N__9297\,
            I => \N__9294\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__9294\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_78\
        );

    \I__1987\ : InMux
    port map (
            O => \N__9291\,
            I => \N__9288\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__9288\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_79\
        );

    \I__1985\ : InMux
    port map (
            O => \N__9285\,
            I => \N__9282\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__9282\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_4\
        );

    \I__1983\ : InMux
    port map (
            O => \N__9279\,
            I => \N__9276\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__9276\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_5\
        );

    \I__1981\ : InMux
    port map (
            O => \N__9273\,
            I => \N__9270\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__9270\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_18\
        );

    \I__1979\ : InMux
    port map (
            O => \N__9267\,
            I => \N__9264\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__9264\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_19\
        );

    \I__1977\ : InMux
    port map (
            O => \N__9261\,
            I => \N__9258\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__9258\,
            I => \N__9255\
        );

    \I__1975\ : Span4Mux_v
    port map (
            O => \N__9255\,
            I => \N__9252\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__9252\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_76\
        );

    \I__1973\ : InMux
    port map (
            O => \N__9249\,
            I => \N__9246\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__9246\,
            I => \N__9243\
        );

    \I__1971\ : Odrv4
    port map (
            O => \N__9243\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_77\
        );

    \I__1970\ : InMux
    port map (
            O => \N__9240\,
            I => \N__9237\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__9237\,
            I => \N__9234\
        );

    \I__1968\ : Odrv4
    port map (
            O => \N__9234\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_39\
        );

    \I__1967\ : InMux
    port map (
            O => \N__9231\,
            I => \N__9228\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__9228\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_3\
        );

    \I__1965\ : InMux
    port map (
            O => \N__9225\,
            I => \N__9222\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__9222\,
            I => \N__9219\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__9219\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_8\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9216\,
            I => \N__9213\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__9213\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_7\
        );

    \I__1960\ : InMux
    port map (
            O => \N__9210\,
            I => \N__9207\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__9207\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_6\
        );

    \I__1958\ : InMux
    port map (
            O => \N__9204\,
            I => \N__9201\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__9201\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_40\
        );

    \I__1956\ : InMux
    port map (
            O => \N__9198\,
            I => \N__9195\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__9195\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_41\
        );

    \I__1954\ : InMux
    port map (
            O => \N__9192\,
            I => \N__9189\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__9189\,
            I => \N__9186\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__9186\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_21\
        );

    \I__1951\ : InMux
    port map (
            O => \N__9183\,
            I => \N__9180\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__9180\,
            I => \N__9177\
        );

    \I__1949\ : Span4Mux_h
    port map (
            O => \N__9177\,
            I => \N__9174\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__9174\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_22\
        );

    \I__1947\ : InMux
    port map (
            O => \N__9171\,
            I => \N__9168\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__9168\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_73\
        );

    \I__1945\ : InMux
    port map (
            O => \N__9165\,
            I => \N__9162\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__9162\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_71\
        );

    \I__1943\ : InMux
    port map (
            O => \N__9159\,
            I => \N__9156\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__9156\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_72\
        );

    \I__1941\ : InMux
    port map (
            O => \N__9153\,
            I => \N__9150\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__9150\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_20\
        );

    \I__1939\ : InMux
    port map (
            O => \N__9147\,
            I => \N__9144\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__9144\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_69\
        );

    \I__1937\ : InMux
    port map (
            O => \N__9141\,
            I => \N__9138\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__9138\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_70\
        );

    \I__1935\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9132\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__9132\,
            I => \N__9129\
        );

    \I__1933\ : Span4Mux_h
    port map (
            O => \N__9129\,
            I => \N__9126\
        );

    \I__1932\ : Odrv4
    port map (
            O => \N__9126\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_15\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__9123\,
            I => \N__9120\
        );

    \I__1930\ : InMux
    port map (
            O => \N__9120\,
            I => \N__9117\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__9117\,
            I => \N__9114\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__9114\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_87\
        );

    \I__1927\ : InMux
    port map (
            O => \N__9111\,
            I => \N__9108\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__9108\,
            I => \N__9105\
        );

    \I__1925\ : Odrv12
    port map (
            O => \N__9105\,
            I => \mosi_1MHz\
        );

    \I__1924\ : CEMux
    port map (
            O => \N__9102\,
            I => \N__9098\
        );

    \I__1923\ : CEMux
    port map (
            O => \N__9101\,
            I => \N__9094\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__9098\,
            I => \N__9091\
        );

    \I__1921\ : InMux
    port map (
            O => \N__9097\,
            I => \N__9085\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__9094\,
            I => \N__9082\
        );

    \I__1919\ : Span4Mux_v
    port map (
            O => \N__9091\,
            I => \N__9073\
        );

    \I__1918\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9068\
        );

    \I__1917\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9068\
        );

    \I__1916\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9064\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__9085\,
            I => \N__9059\
        );

    \I__1914\ : Span4Mux_h
    port map (
            O => \N__9082\,
            I => \N__9059\
        );

    \I__1913\ : InMux
    port map (
            O => \N__9081\,
            I => \N__9056\
        );

    \I__1912\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9047\
        );

    \I__1911\ : InMux
    port map (
            O => \N__9079\,
            I => \N__9047\
        );

    \I__1910\ : InMux
    port map (
            O => \N__9078\,
            I => \N__9047\
        );

    \I__1909\ : InMux
    port map (
            O => \N__9077\,
            I => \N__9047\
        );

    \I__1908\ : InMux
    port map (
            O => \N__9076\,
            I => \N__9044\
        );

    \I__1907\ : Span4Mux_h
    port map (
            O => \N__9073\,
            I => \N__9039\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__9068\,
            I => \N__9039\
        );

    \I__1905\ : InMux
    port map (
            O => \N__9067\,
            I => \N__9036\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__9064\,
            I => \counter_RNISR1F_2\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__9059\,
            I => \counter_RNISR1F_2\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__9056\,
            I => \counter_RNISR1F_2\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__9047\,
            I => \counter_RNISR1F_2\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__9044\,
            I => \counter_RNISR1F_2\
        );

    \I__1899\ : Odrv4
    port map (
            O => \N__9039\,
            I => \counter_RNISR1F_2\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__9036\,
            I => \counter_RNISR1F_2\
        );

    \I__1897\ : InMux
    port map (
            O => \N__9021\,
            I => \N__9018\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__9018\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_85\
        );

    \I__1895\ : InMux
    port map (
            O => \N__9015\,
            I => \N__9012\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__9012\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_82\
        );

    \I__1893\ : InMux
    port map (
            O => \N__9009\,
            I => \N__9006\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__9006\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_83\
        );

    \I__1891\ : InMux
    port map (
            O => \N__9003\,
            I => \N__9000\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__9000\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_84\
        );

    \I__1889\ : InMux
    port map (
            O => \N__8997\,
            I => \N__8994\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8994\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_16\
        );

    \I__1887\ : InMux
    port map (
            O => \N__8991\,
            I => \N__8988\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__8988\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_80\
        );

    \I__1885\ : InMux
    port map (
            O => \N__8985\,
            I => \N__8982\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__8982\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_74\
        );

    \I__1883\ : InMux
    port map (
            O => \N__8979\,
            I => \N__8976\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__8976\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_75\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8973\,
            I => \N__8970\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__8970\,
            I => \N__8967\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__8967\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_67\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8964\,
            I => \N__8961\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8961\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_42\
        );

    \I__1876\ : InMux
    port map (
            O => \N__8958\,
            I => \N__8955\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8955\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_43\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8952\,
            I => \N__8949\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__8949\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_44\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8946\,
            I => \N__8943\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8943\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_45\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8940\,
            I => \N__8937\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__8937\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_46\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8934\,
            I => \N__8931\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8931\,
            I => \N__8928\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__8928\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_47\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8925\,
            I => \N__8922\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8922\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_68\
        );

    \I__1863\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8916\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__8916\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_48\
        );

    \I__1861\ : InMux
    port map (
            O => \N__8913\,
            I => \N__8910\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__8910\,
            I => \N__8907\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__8907\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_15\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8901\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__8901\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_50\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8898\,
            I => \N__8895\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__8895\,
            I => \N__8892\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__8892\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_51\
        );

    \I__1853\ : InMux
    port map (
            O => \N__8889\,
            I => \N__8886\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__8886\,
            I => \N__8883\
        );

    \I__1851\ : Odrv4
    port map (
            O => \N__8883\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_33\
        );

    \I__1850\ : InMux
    port map (
            O => \N__8880\,
            I => \N__8877\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__8877\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_34\
        );

    \I__1848\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8871\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__8871\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_66\
        );

    \I__1846\ : InMux
    port map (
            O => \N__8868\,
            I => \N__8865\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__8865\,
            I => \N__8862\
        );

    \I__1844\ : Odrv4
    port map (
            O => \N__8862\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_64\
        );

    \I__1843\ : InMux
    port map (
            O => \N__8859\,
            I => \N__8856\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__8856\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_65\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8853\,
            I => \N__8850\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8850\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_13\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8844\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8844\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_14\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8837\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8840\,
            I => \N__8834\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8837\,
            I => \N__8831\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__8834\,
            I => \N__8828\
        );

    \I__1833\ : Span4Mux_h
    port map (
            O => \N__8831\,
            I => \N__8825\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__8828\,
            I => \switch_clk_1MHz_inst_delay_inst_delay_reg_15\
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__8825\,
            I => \switch_clk_1MHz_inst_delay_inst_delay_reg_15\
        );

    \I__1830\ : InMux
    port map (
            O => \N__8820\,
            I => \N__8817\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__8817\,
            I => \N__8813\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8810\
        );

    \I__1827\ : Odrv4
    port map (
            O => \N__8813\,
            I => \config_register_latched_dec_inst.STATCNF_1Z0Z_0\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__8810\,
            I => \config_register_latched_dec_inst.STATCNF_1Z0Z_0\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8805\,
            I => \N__8801\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__8804\,
            I => \N__8798\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8801\,
            I => \N__8795\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8798\,
            I => \N__8792\
        );

    \I__1821\ : Span4Mux_h
    port map (
            O => \N__8795\,
            I => \N__8786\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8792\,
            I => \N__8786\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__8791\,
            I => \N__8783\
        );

    \I__1818\ : Span4Mux_h
    port map (
            O => \N__8786\,
            I => \N__8778\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8783\,
            I => \N__8773\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8782\,
            I => \N__8773\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8781\,
            I => \N__8770\
        );

    \I__1814\ : Span4Mux_v
    port map (
            O => \N__8778\,
            I => \N__8767\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8773\,
            I => \N__8764\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8770\,
            I => \N__8761\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__8767\,
            I => \N__8758\
        );

    \I__1810\ : Sp12to4
    port map (
            O => \N__8764\,
            I => \N__8755\
        );

    \I__1809\ : Sp12to4
    port map (
            O => \N__8761\,
            I => \N__8752\
        );

    \I__1808\ : Sp12to4
    port map (
            O => \N__8758\,
            I => \N__8747\
        );

    \I__1807\ : Span12Mux_v
    port map (
            O => \N__8755\,
            I => \N__8747\
        );

    \I__1806\ : Span12Mux_v
    port map (
            O => \N__8752\,
            I => \N__8744\
        );

    \I__1805\ : Odrv12
    port map (
            O => \N__8747\,
            I => \RST_N_c\
        );

    \I__1804\ : Odrv12
    port map (
            O => \N__8744\,
            I => \RST_N_c\
        );

    \I__1803\ : IoInMux
    port map (
            O => \N__8739\,
            I => \N__8736\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8736\,
            I => \N__8733\
        );

    \I__1801\ : IoSpan4Mux
    port map (
            O => \N__8733\,
            I => \N__8730\
        );

    \I__1800\ : Span4Mux_s3_h
    port map (
            O => \N__8730\,
            I => \N__8727\
        );

    \I__1799\ : Sp12to4
    port map (
            O => \N__8727\,
            I => \N__8723\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__8726\,
            I => \N__8720\
        );

    \I__1797\ : Span12Mux_h
    port map (
            O => \N__8723\,
            I => \N__8717\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8720\,
            I => \N__8714\
        );

    \I__1795\ : Span12Mux_h
    port map (
            O => \N__8717\,
            I => \N__8711\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__8714\,
            I => \N__8708\
        );

    \I__1793\ : Span12Mux_v
    port map (
            O => \N__8711\,
            I => \N__8700\
        );

    \I__1792\ : Span4Mux_v
    port map (
            O => \N__8708\,
            I => \N__8697\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8707\,
            I => \N__8694\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8706\,
            I => \N__8689\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8705\,
            I => \N__8689\
        );

    \I__1788\ : InMux
    port map (
            O => \N__8704\,
            I => \N__8684\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8703\,
            I => \N__8684\
        );

    \I__1786\ : Odrv12
    port map (
            O => \N__8700\,
            I => sel_output_c
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__8697\,
            I => sel_output_c
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8694\,
            I => sel_output_c
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8689\,
            I => sel_output_c
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8684\,
            I => sel_output_c
        );

    \I__1781\ : InMux
    port map (
            O => \N__8673\,
            I => \N__8670\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8670\,
            I => \N__8667\
        );

    \I__1779\ : Span4Mux_v
    port map (
            O => \N__8667\,
            I => \N__8662\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8659\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8665\,
            I => \N__8656\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__8662\,
            I => \config_register_latched_dec_inst.STATSRZ0Z_0\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__8659\,
            I => \config_register_latched_dec_inst.STATSRZ0Z_0\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__8656\,
            I => \config_register_latched_dec_inst.STATSRZ0Z_0\
        );

    \I__1773\ : InMux
    port map (
            O => \N__8649\,
            I => \N__8646\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8646\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_81\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8643\,
            I => \N__8640\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8640\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_86\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8637\,
            I => \N__8634\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8634\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_49\
        );

    \I__1767\ : InMux
    port map (
            O => \N__8631\,
            I => \N__8628\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__8628\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_13\
        );

    \I__1765\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8622\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8622\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_14\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8616\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__8616\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_52\
        );

    \I__1761\ : InMux
    port map (
            O => \N__8613\,
            I => \N__8610\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__8610\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_53\
        );

    \I__1759\ : InMux
    port map (
            O => \N__8607\,
            I => \N__8604\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__8604\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_11\
        );

    \I__1757\ : InMux
    port map (
            O => \N__8601\,
            I => \N__8598\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8598\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_9\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8592\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__8592\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_10\
        );

    \I__1753\ : InMux
    port map (
            O => \N__8589\,
            I => \N__8586\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__8586\,
            I => \N__8583\
        );

    \I__1751\ : Odrv4
    port map (
            O => \N__8583\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_8\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8580\,
            I => \N__8577\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__8577\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_9\
        );

    \I__1748\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8571\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__8571\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_10\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8565\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__8565\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_11\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8559\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8559\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_12\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__8556\,
            I => \N__8552\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8555\,
            I => \N__8546\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8546\
        );

    \I__1739\ : InMux
    port map (
            O => \N__8551\,
            I => \N__8543\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__8546\,
            I => \N__8540\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__8543\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_0\
        );

    \I__1736\ : Odrv4
    port map (
            O => \N__8540\,
            I => \config_register_latched_dec_inst.DYNSRZ0Z_0\
        );

    \I__1735\ : InMux
    port map (
            O => \N__8535\,
            I => \N__8529\
        );

    \I__1734\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8529\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8529\,
            I => \N__8526\
        );

    \I__1732\ : Span12Mux_h
    port map (
            O => \N__8526\,
            I => \N__8523\
        );

    \I__1731\ : Span12Mux_h
    port map (
            O => \N__8523\,
            I => \N__8520\
        );

    \I__1730\ : Odrv12
    port map (
            O => \N__8520\,
            I => miso_input_c
        );

    \I__1729\ : CEMux
    port map (
            O => \N__8517\,
            I => \N__8514\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__8514\,
            I => \N__8511\
        );

    \I__1727\ : Span4Mux_h
    port map (
            O => \N__8511\,
            I => \N__8508\
        );

    \I__1726\ : Odrv4
    port map (
            O => \N__8508\,
            I => \delay_reg_RNI7S8U1_15\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8505\,
            I => \N__8502\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__8502\,
            I => \N__8499\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__8499\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_32\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8493\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__8493\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_54\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8490\,
            I => \N__8487\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8487\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_12\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8484\,
            I => \N__8481\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8481\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_4\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8478\,
            I => \N__8475\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8475\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_7\
        );

    \I__1714\ : InMux
    port map (
            O => \N__8472\,
            I => \N__8469\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__8469\,
            I => \N__8466\
        );

    \I__1712\ : Span4Mux_h
    port map (
            O => \N__8466\,
            I => \N__8463\
        );

    \I__1711\ : Odrv4
    port map (
            O => \N__8463\,
            I => \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_2\
        );

    \I__1710\ : InMux
    port map (
            O => \N__8460\,
            I => \N__8454\
        );

    \I__1709\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8451\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8458\,
            I => \N__8446\
        );

    \I__1707\ : InMux
    port map (
            O => \N__8457\,
            I => \N__8446\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8454\,
            I => \N_4_0\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__8451\,
            I => \N_4_0\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__8446\,
            I => \N_4_0\
        );

    \I__1703\ : IoInMux
    port map (
            O => \N__8439\,
            I => \N__8436\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__8436\,
            I => \N__8433\
        );

    \I__1701\ : Span4Mux_s3_v
    port map (
            O => \N__8433\,
            I => \N__8430\
        );

    \I__1700\ : Span4Mux_h
    port map (
            O => \N__8430\,
            I => \N__8427\
        );

    \I__1699\ : Sp12to4
    port map (
            O => \N__8427\,
            I => \N__8424\
        );

    \I__1698\ : Span12Mux_v
    port map (
            O => \N__8424\,
            I => \N__8421\
        );

    \I__1697\ : Span12Mux_h
    port map (
            O => \N__8421\,
            I => \N__8417\
        );

    \I__1696\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8414\
        );

    \I__1695\ : Odrv12
    port map (
            O => \N__8417\,
            I => clk_output_c
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__8414\,
            I => clk_output_c
        );

    \I__1693\ : InMux
    port map (
            O => \N__8409\,
            I => \N__8405\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8402\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__8405\,
            I => \switch_clk_2MHz_inst_delay_inst_delay_reg_6\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__8402\,
            I => \switch_clk_2MHz_inst_delay_inst_delay_reg_6\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8397\,
            I => \N__8394\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__8394\,
            I => \N__8391\
        );

    \I__1687\ : Odrv4
    port map (
            O => \N__8391\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_2\
        );

    \I__1686\ : InMux
    port map (
            O => \N__8388\,
            I => \N__8385\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__8385\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_3\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8382\,
            I => \N__8379\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8379\,
            I => \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_3\
        );

    \I__1682\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8373\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__8373\,
            I => \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_4\
        );

    \I__1680\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8367\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8367\,
            I => \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_5\
        );

    \I__1678\ : CEMux
    port map (
            O => \N__8364\,
            I => \N__8361\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__8361\,
            I => \N__8358\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__8358\,
            I => \config_register_latched_dec_inst.N_381_i_i\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8355\,
            I => \N__8352\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8352\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_55\
        );

    \I__1673\ : InMux
    port map (
            O => \N__8349\,
            I => \N__8346\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8346\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_56\
        );

    \I__1671\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8340\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__8340\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_62\
        );

    \I__1669\ : InMux
    port map (
            O => \N__8337\,
            I => \N__8334\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__8334\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_63\
        );

    \I__1667\ : InMux
    port map (
            O => \N__8331\,
            I => \N__8328\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__8328\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_31\
        );

    \I__1665\ : InMux
    port map (
            O => \N__8325\,
            I => \N__8322\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__8322\,
            I => \N__8319\
        );

    \I__1663\ : Odrv4
    port map (
            O => \N__8319\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1662\ : CascadeMux
    port map (
            O => \N__8316\,
            I => \N__8309\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__8315\,
            I => \N__8306\
        );

    \I__1660\ : InMux
    port map (
            O => \N__8314\,
            I => \N__8302\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8313\,
            I => \N__8297\
        );

    \I__1658\ : InMux
    port map (
            O => \N__8312\,
            I => \N__8297\
        );

    \I__1657\ : InMux
    port map (
            O => \N__8309\,
            I => \N__8292\
        );

    \I__1656\ : InMux
    port map (
            O => \N__8306\,
            I => \N__8292\
        );

    \I__1655\ : InMux
    port map (
            O => \N__8305\,
            I => \N__8289\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__8302\,
            I => divisor_inst_counter_1
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__8297\,
            I => divisor_inst_counter_1
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__8292\,
            I => divisor_inst_counter_1
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__8289\,
            I => divisor_inst_counter_1
        );

    \I__1650\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8269\
        );

    \I__1649\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8269\
        );

    \I__1648\ : InMux
    port map (
            O => \N__8278\,
            I => \N__8260\
        );

    \I__1647\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8260\
        );

    \I__1646\ : InMux
    port map (
            O => \N__8276\,
            I => \N__8260\
        );

    \I__1645\ : InMux
    port map (
            O => \N__8275\,
            I => \N__8260\
        );

    \I__1644\ : InMux
    port map (
            O => \N__8274\,
            I => \N__8257\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__8269\,
            I => divisor_inst_counter_0
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__8260\,
            I => divisor_inst_counter_0
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__8257\,
            I => divisor_inst_counter_0
        );

    \I__1640\ : InMux
    port map (
            O => \N__8250\,
            I => \N__8247\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__8247\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_reg_0_6\
        );

    \I__1638\ : InMux
    port map (
            O => \N__8244\,
            I => \N__8241\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__8241\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_5\
        );

    \I__1636\ : InMux
    port map (
            O => \N__8238\,
            I => \N__8227\
        );

    \I__1635\ : InMux
    port map (
            O => \N__8237\,
            I => \N__8227\
        );

    \I__1634\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8227\
        );

    \I__1633\ : InMux
    port map (
            O => \N__8235\,
            I => \N__8224\
        );

    \I__1632\ : InMux
    port map (
            O => \N__8234\,
            I => \N__8221\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__8227\,
            I => \divisor_inst_2.counterZ0Z_0\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__8224\,
            I => \divisor_inst_2.counterZ0Z_0\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__8221\,
            I => \divisor_inst_2.counterZ0Z_0\
        );

    \I__1628\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8207\
        );

    \I__1627\ : InMux
    port map (
            O => \N__8213\,
            I => \N__8207\
        );

    \I__1626\ : InMux
    port map (
            O => \N__8212\,
            I => \N__8204\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__8207\,
            I => \divisor_inst_2.counterZ0Z_2\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__8204\,
            I => \divisor_inst_2.counterZ0Z_2\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__8199\,
            I => \N__8195\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__8198\,
            I => \N__8190\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8195\,
            I => \N__8183\
        );

    \I__1620\ : InMux
    port map (
            O => \N__8194\,
            I => \N__8183\
        );

    \I__1619\ : InMux
    port map (
            O => \N__8193\,
            I => \N__8183\
        );

    \I__1618\ : InMux
    port map (
            O => \N__8190\,
            I => \N__8180\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__8183\,
            I => \divisor_inst_2.counterZ0Z_1\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__8180\,
            I => \divisor_inst_2.counterZ0Z_1\
        );

    \I__1615\ : InMux
    port map (
            O => \N__8175\,
            I => \N__8172\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__8172\,
            I => \switch_clk_2MHz_inst.SEL_0_RNI98MZ0Z31\
        );

    \I__1613\ : InMux
    port map (
            O => \N__8169\,
            I => \N__8165\
        );

    \I__1612\ : InMux
    port map (
            O => \N__8168\,
            I => \N__8162\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__8165\,
            I => \N_3_0\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__8162\,
            I => \N_3_0\
        );

    \I__1609\ : InMux
    port map (
            O => \N__8157\,
            I => \N__8151\
        );

    \I__1608\ : InMux
    port map (
            O => \N__8156\,
            I => \N__8148\
        );

    \I__1607\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8143\
        );

    \I__1606\ : InMux
    port map (
            O => \N__8154\,
            I => \N__8143\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__8151\,
            I => flag_signal
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__8148\,
            I => flag_signal
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__8143\,
            I => flag_signal
        );

    \I__1602\ : InMux
    port map (
            O => \N__8136\,
            I => \N__8133\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__8133\,
            I => \N__8130\
        );

    \I__1600\ : Odrv4
    port map (
            O => \N__8130\,
            I => \switch_clk_1MHz_inst.flag_input_regZ0\
        );

    \I__1599\ : InMux
    port map (
            O => \N__8127\,
            I => \N__8122\
        );

    \I__1598\ : InMux
    port map (
            O => \N__8126\,
            I => \N__8119\
        );

    \I__1597\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8116\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__8122\,
            I => \clk_continuous_1MHz\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__8119\,
            I => \clk_continuous_1MHz\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__8116\,
            I => \clk_continuous_1MHz\
        );

    \I__1593\ : InMux
    port map (
            O => \N__8109\,
            I => \N__8106\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__8106\,
            I => \N__8103\
        );

    \I__1591\ : Odrv4
    port map (
            O => \N__8103\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_1\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__8100\,
            I => \N__8097\
        );

    \I__1589\ : InMux
    port map (
            O => \N__8097\,
            I => \N__8094\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__8094\,
            I => \N__8091\
        );

    \I__1587\ : Odrv4
    port map (
            O => \N__8091\,
            I => \switch_clk_1MHz_inst.N_91_0\
        );

    \I__1586\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8085\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__8085\,
            I => \N__8078\
        );

    \I__1584\ : InMux
    port map (
            O => \N__8084\,
            I => \N__8071\
        );

    \I__1583\ : InMux
    port map (
            O => \N__8083\,
            I => \N__8071\
        );

    \I__1582\ : InMux
    port map (
            O => \N__8082\,
            I => \N__8071\
        );

    \I__1581\ : InMux
    port map (
            O => \N__8081\,
            I => \N__8068\
        );

    \I__1580\ : Odrv4
    port map (
            O => \N__8078\,
            I => \switch_clk_1MHz_inst.N_90_li\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__8071\,
            I => \switch_clk_1MHz_inst.N_90_li\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__8068\,
            I => \switch_clk_1MHz_inst.N_90_li\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__8061\,
            I => \N__8057\
        );

    \I__1576\ : InMux
    port map (
            O => \N__8060\,
            I => \N__8053\
        );

    \I__1575\ : InMux
    port map (
            O => \N__8057\,
            I => \N__8048\
        );

    \I__1574\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8048\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__8053\,
            I => \switch_clk_1MHz_inst.counter_dinZ0Z_3\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__8048\,
            I => \switch_clk_1MHz_inst.counter_dinZ0Z_3\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__8043\,
            I => \N__8039\
        );

    \I__1570\ : InMux
    port map (
            O => \N__8042\,
            I => \N__8034\
        );

    \I__1569\ : InMux
    port map (
            O => \N__8039\,
            I => \N__8034\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__8034\,
            I => \switch_clk_1MHz_inst.CLK_uCZ0\
        );

    \I__1567\ : InMux
    port map (
            O => \N__8031\,
            I => \N__8028\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__8028\,
            I => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_0\
        );

    \I__1565\ : InMux
    port map (
            O => \N__8025\,
            I => \N__8021\
        );

    \I__1564\ : InMux
    port map (
            O => \N__8024\,
            I => \N__8018\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__8021\,
            I => \aux_selection_1MHz_0\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__8018\,
            I => \aux_selection_1MHz_0\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__8013\,
            I => \N_4_0_cascade_\
        );

    \I__1560\ : InMux
    port map (
            O => \N__8010\,
            I => \N__8007\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__8007\,
            I => \N__8004\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__8004\,
            I => \config_register_latched_dec_inst.STATCNF_1_RNO_0Z0Z_0\
        );

    \I__1557\ : InMux
    port map (
            O => \N__8001\,
            I => \N__7998\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7998\,
            I => \N_2_0\
        );

    \I__1555\ : InMux
    port map (
            O => \N__7995\,
            I => \N__7959\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7994\,
            I => \N__7959\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7993\,
            I => \N__7959\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7992\,
            I => \N__7959\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7991\,
            I => \N__7959\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7990\,
            I => \N__7956\
        );

    \I__1549\ : InMux
    port map (
            O => \N__7989\,
            I => \N__7943\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7988\,
            I => \N__7943\
        );

    \I__1547\ : InMux
    port map (
            O => \N__7987\,
            I => \N__7943\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7986\,
            I => \N__7943\
        );

    \I__1545\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7943\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7943\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7983\,
            I => \N__7934\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7982\,
            I => \N__7934\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7981\,
            I => \N__7934\
        );

    \I__1540\ : InMux
    port map (
            O => \N__7980\,
            I => \N__7934\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7979\,
            I => \N__7921\
        );

    \I__1538\ : InMux
    port map (
            O => \N__7978\,
            I => \N__7921\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7977\,
            I => \N__7921\
        );

    \I__1536\ : InMux
    port map (
            O => \N__7976\,
            I => \N__7921\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7975\,
            I => \N__7921\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7974\,
            I => \N__7921\
        );

    \I__1533\ : CascadeMux
    port map (
            O => \N__7973\,
            I => \N__7904\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__7972\,
            I => \N__7901\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__7971\,
            I => \N__7898\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__7970\,
            I => \N__7895\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__7959\,
            I => \N__7851\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7956\,
            I => \N__7851\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7943\,
            I => \N__7851\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__7934\,
            I => \N__7851\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__7921\,
            I => \N__7848\
        );

    \I__1524\ : InMux
    port map (
            O => \N__7920\,
            I => \N__7833\
        );

    \I__1523\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7833\
        );

    \I__1522\ : InMux
    port map (
            O => \N__7918\,
            I => \N__7833\
        );

    \I__1521\ : InMux
    port map (
            O => \N__7917\,
            I => \N__7833\
        );

    \I__1520\ : InMux
    port map (
            O => \N__7916\,
            I => \N__7833\
        );

    \I__1519\ : InMux
    port map (
            O => \N__7915\,
            I => \N__7833\
        );

    \I__1518\ : InMux
    port map (
            O => \N__7914\,
            I => \N__7833\
        );

    \I__1517\ : InMux
    port map (
            O => \N__7913\,
            I => \N__7797\
        );

    \I__1516\ : InMux
    port map (
            O => \N__7912\,
            I => \N__7797\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7911\,
            I => \N__7797\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7797\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7797\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7792\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7907\,
            I => \N__7792\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7904\,
            I => \N__7781\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7901\,
            I => \N__7781\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7898\,
            I => \N__7781\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7895\,
            I => \N__7781\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7894\,
            I => \N__7781\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7893\,
            I => \N__7764\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7892\,
            I => \N__7764\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7891\,
            I => \N__7764\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7890\,
            I => \N__7764\
        );

    \I__1501\ : InMux
    port map (
            O => \N__7889\,
            I => \N__7764\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7888\,
            I => \N__7764\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7887\,
            I => \N__7764\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7886\,
            I => \N__7764\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7885\,
            I => \N__7753\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7884\,
            I => \N__7753\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7883\,
            I => \N__7753\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7882\,
            I => \N__7753\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7753\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7738\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7879\,
            I => \N__7738\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7738\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7738\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7738\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7738\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7874\,
            I => \N__7738\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7873\,
            I => \N__7721\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7872\,
            I => \N__7721\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7871\,
            I => \N__7721\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7870\,
            I => \N__7721\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7869\,
            I => \N__7721\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7868\,
            I => \N__7721\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7867\,
            I => \N__7721\
        );

    \I__1478\ : InMux
    port map (
            O => \N__7866\,
            I => \N__7721\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7865\,
            I => \N__7708\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7864\,
            I => \N__7708\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7863\,
            I => \N__7708\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7862\,
            I => \N__7708\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7861\,
            I => \N__7708\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7860\,
            I => \N__7708\
        );

    \I__1471\ : Span4Mux_v
    port map (
            O => \N__7851\,
            I => \N__7699\
        );

    \I__1470\ : Span4Mux_v
    port map (
            O => \N__7848\,
            I => \N__7699\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7833\,
            I => \N__7699\
        );

    \I__1468\ : InMux
    port map (
            O => \N__7832\,
            I => \N__7696\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7831\,
            I => \N__7685\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7830\,
            I => \N__7682\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7829\,
            I => \N__7665\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7828\,
            I => \N__7665\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7827\,
            I => \N__7665\
        );

    \I__1462\ : InMux
    port map (
            O => \N__7826\,
            I => \N__7665\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7825\,
            I => \N__7665\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7824\,
            I => \N__7665\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7665\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7822\,
            I => \N__7665\
        );

    \I__1457\ : InMux
    port map (
            O => \N__7821\,
            I => \N__7648\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7820\,
            I => \N__7648\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7819\,
            I => \N__7648\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7818\,
            I => \N__7648\
        );

    \I__1453\ : InMux
    port map (
            O => \N__7817\,
            I => \N__7648\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7816\,
            I => \N__7648\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7815\,
            I => \N__7648\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7814\,
            I => \N__7648\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7813\,
            I => \N__7637\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7637\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7637\
        );

    \I__1446\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7637\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7637\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7808\,
            I => \N__7634\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7797\,
            I => \N__7631\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__7792\,
            I => \N__7622\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7781\,
            I => \N__7622\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__7764\,
            I => \N__7622\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__7753\,
            I => \N__7622\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__7738\,
            I => \N__7613\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__7721\,
            I => \N__7613\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7708\,
            I => \N__7613\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7707\,
            I => \N__7600\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7706\,
            I => \N__7600\
        );

    \I__1433\ : Span4Mux_h
    port map (
            O => \N__7699\,
            I => \N__7595\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7696\,
            I => \N__7595\
        );

    \I__1431\ : InMux
    port map (
            O => \N__7695\,
            I => \N__7584\
        );

    \I__1430\ : InMux
    port map (
            O => \N__7694\,
            I => \N__7584\
        );

    \I__1429\ : InMux
    port map (
            O => \N__7693\,
            I => \N__7584\
        );

    \I__1428\ : InMux
    port map (
            O => \N__7692\,
            I => \N__7584\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7691\,
            I => \N__7575\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7690\,
            I => \N__7575\
        );

    \I__1425\ : InMux
    port map (
            O => \N__7689\,
            I => \N__7575\
        );

    \I__1424\ : InMux
    port map (
            O => \N__7688\,
            I => \N__7575\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__7685\,
            I => \N__7572\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7682\,
            I => \N__7563\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__7665\,
            I => \N__7563\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__7648\,
            I => \N__7563\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__7637\,
            I => \N__7563\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__7634\,
            I => \N__7556\
        );

    \I__1417\ : Span4Mux_s2_h
    port map (
            O => \N__7631\,
            I => \N__7556\
        );

    \I__1416\ : Span4Mux_v
    port map (
            O => \N__7622\,
            I => \N__7556\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7621\,
            I => \N__7551\
        );

    \I__1414\ : InMux
    port map (
            O => \N__7620\,
            I => \N__7551\
        );

    \I__1413\ : Span4Mux_h
    port map (
            O => \N__7613\,
            I => \N__7548\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7537\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7611\,
            I => \N__7537\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7610\,
            I => \N__7537\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7609\,
            I => \N__7537\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7608\,
            I => \N__7537\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7607\,
            I => \N__7532\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7606\,
            I => \N__7532\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7605\,
            I => \N__7529\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7600\,
            I => \N__7524\
        );

    \I__1403\ : Span4Mux_v
    port map (
            O => \N__7595\,
            I => \N__7524\
        );

    \I__1402\ : InMux
    port map (
            O => \N__7594\,
            I => \N__7519\
        );

    \I__1401\ : InMux
    port map (
            O => \N__7593\,
            I => \N__7519\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7584\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_0\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7575\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_0\
        );

    \I__1398\ : Odrv4
    port map (
            O => \N__7572\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_0\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__7563\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_0\
        );

    \I__1396\ : Odrv4
    port map (
            O => \N__7556\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_0\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__7551\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_0\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__7548\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_0\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7537\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_0\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7532\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_0\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7529\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_0\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__7524\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_0\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__7519\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_0\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__7494\,
            I => \N__7491\
        );

    \I__1387\ : InMux
    port map (
            O => \N__7491\,
            I => \N__7484\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__7490\,
            I => \N__7481\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__7489\,
            I => \N__7477\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7488\,
            I => \N__7472\
        );

    \I__1383\ : InMux
    port map (
            O => \N__7487\,
            I => \N__7472\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__7484\,
            I => \N__7469\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7481\,
            I => \N__7466\
        );

    \I__1380\ : InMux
    port map (
            O => \N__7480\,
            I => \N__7457\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7477\,
            I => \N__7457\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__7472\,
            I => \N__7454\
        );

    \I__1377\ : Span4Mux_v
    port map (
            O => \N__7469\,
            I => \N__7449\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__7466\,
            I => \N__7449\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7465\,
            I => \N__7446\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7464\,
            I => \N__7443\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7463\,
            I => \N__7438\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7462\,
            I => \N__7438\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7457\,
            I => \N__7433\
        );

    \I__1370\ : Span4Mux_h
    port map (
            O => \N__7454\,
            I => \N__7433\
        );

    \I__1369\ : Span4Mux_v
    port map (
            O => \N__7449\,
            I => \N__7430\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7446\,
            I => \switch_clk_2MHz_inst.current_state_fast_1_repZ0Z1\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__7443\,
            I => \switch_clk_2MHz_inst.current_state_fast_1_repZ0Z1\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__7438\,
            I => \switch_clk_2MHz_inst.current_state_fast_1_repZ0Z1\
        );

    \I__1365\ : Odrv4
    port map (
            O => \N__7433\,
            I => \switch_clk_2MHz_inst.current_state_fast_1_repZ0Z1\
        );

    \I__1364\ : Odrv4
    port map (
            O => \N__7430\,
            I => \switch_clk_2MHz_inst.current_state_fast_1_repZ0Z1\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7419\,
            I => \N__7412\
        );

    \I__1362\ : CascadeMux
    port map (
            O => \N__7418\,
            I => \N__7408\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7417\,
            I => \N__7394\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7416\,
            I => \N__7394\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7415\,
            I => \N__7391\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__7412\,
            I => \N__7388\
        );

    \I__1357\ : InMux
    port map (
            O => \N__7411\,
            I => \N__7381\
        );

    \I__1356\ : InMux
    port map (
            O => \N__7408\,
            I => \N__7376\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7407\,
            I => \N__7376\
        );

    \I__1354\ : InMux
    port map (
            O => \N__7406\,
            I => \N__7367\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7405\,
            I => \N__7367\
        );

    \I__1352\ : InMux
    port map (
            O => \N__7404\,
            I => \N__7367\
        );

    \I__1351\ : InMux
    port map (
            O => \N__7403\,
            I => \N__7367\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7402\,
            I => \N__7364\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7401\,
            I => \N__7357\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7400\,
            I => \N__7357\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7399\,
            I => \N__7357\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__7394\,
            I => \N__7354\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__7391\,
            I => \N__7349\
        );

    \I__1344\ : Span4Mux_h
    port map (
            O => \N__7388\,
            I => \N__7349\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7387\,
            I => \N__7344\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7344\
        );

    \I__1341\ : CEMux
    port map (
            O => \N__7385\,
            I => \N__7339\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7384\,
            I => \N__7339\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__7381\,
            I => \N__7334\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__7376\,
            I => \N__7334\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__7367\,
            I => \clk_out_RNI3LEM\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7364\,
            I => \clk_out_RNI3LEM\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__7357\,
            I => \clk_out_RNI3LEM\
        );

    \I__1334\ : Odrv12
    port map (
            O => \N__7354\,
            I => \clk_out_RNI3LEM\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__7349\,
            I => \clk_out_RNI3LEM\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__7344\,
            I => \clk_out_RNI3LEM\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__7339\,
            I => \clk_out_RNI3LEM\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__7334\,
            I => \clk_out_RNI3LEM\
        );

    \I__1329\ : InMux
    port map (
            O => \N__7317\,
            I => \N__7314\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__7314\,
            I => \switch_clk_2MHz_inst.SEL_0_RNIC97QZ0Z_0\
        );

    \I__1327\ : CascadeMux
    port map (
            O => \N__7311\,
            I => \switch_clk_2MHz_inst.SEL_0_RNIC97QZ0Z_0_cascade_\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7308\,
            I => \N__7305\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__7305\,
            I => \switch_clk_2MHz_inst.SEL_0_RNIC97QZ0\
        );

    \I__1324\ : CascadeMux
    port map (
            O => \N__7302\,
            I => \switch_clk_2MHz_inst.N_91_li_cascade_\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7299\,
            I => \N__7296\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__7296\,
            I => \N__7293\
        );

    \I__1321\ : Span4Mux_h
    port map (
            O => \N__7293\,
            I => \N__7285\
        );

    \I__1320\ : InMux
    port map (
            O => \N__7292\,
            I => \N__7276\
        );

    \I__1319\ : InMux
    port map (
            O => \N__7291\,
            I => \N__7276\
        );

    \I__1318\ : InMux
    port map (
            O => \N__7290\,
            I => \N__7276\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7289\,
            I => \N__7276\
        );

    \I__1316\ : InMux
    port map (
            O => \N__7288\,
            I => \N__7273\
        );

    \I__1315\ : Odrv4
    port map (
            O => \N__7285\,
            I => \clk_continuous_2MHz\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__7276\,
            I => \clk_continuous_2MHz\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__7273\,
            I => \clk_continuous_2MHz\
        );

    \I__1312\ : IoInMux
    port map (
            O => \N__7266\,
            I => \N__7263\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__7263\,
            I => \N__7260\
        );

    \I__1310\ : Span4Mux_s2_h
    port map (
            O => \N__7260\,
            I => \N__7257\
        );

    \I__1309\ : Span4Mux_v
    port map (
            O => \N__7257\,
            I => \N__7254\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__7254\,
            I => \switch_clk_2MHz_inst.current_state_fast_fast_RNI0KTVZ0Z_1\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__7251\,
            I => \N__7248\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7248\,
            I => \N__7243\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__7247\,
            I => \N__7240\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__7246\,
            I => \N__7236\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__7243\,
            I => \N__7232\
        );

    \I__1302\ : InMux
    port map (
            O => \N__7240\,
            I => \N__7229\
        );

    \I__1301\ : InMux
    port map (
            O => \N__7239\,
            I => \N__7222\
        );

    \I__1300\ : InMux
    port map (
            O => \N__7236\,
            I => \N__7222\
        );

    \I__1299\ : InMux
    port map (
            O => \N__7235\,
            I => \N__7222\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__7232\,
            I => \switch_clk_2MHz_inst.N_114_0\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__7229\,
            I => \switch_clk_2MHz_inst.N_114_0\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__7222\,
            I => \switch_clk_2MHz_inst.N_114_0\
        );

    \I__1295\ : InMux
    port map (
            O => \N__7215\,
            I => \N__7211\
        );

    \I__1294\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7208\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__7211\,
            I => \switch_clk_2MHz_inst.current_state_fast_fastZ0Z_1\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__7208\,
            I => \switch_clk_2MHz_inst.current_state_fast_fastZ0Z_1\
        );

    \I__1291\ : InMux
    port map (
            O => \N__7203\,
            I => \N__7200\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__7200\,
            I => \mosi_2MHz\
        );

    \I__1289\ : IoInMux
    port map (
            O => \N__7197\,
            I => \N__7194\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__7194\,
            I => \N__7191\
        );

    \I__1287\ : Span4Mux_s2_h
    port map (
            O => \N__7191\,
            I => \N__7188\
        );

    \I__1286\ : Sp12to4
    port map (
            O => \N__7188\,
            I => \N__7185\
        );

    \I__1285\ : Span12Mux_s10_v
    port map (
            O => \N__7185\,
            I => \N__7182\
        );

    \I__1284\ : Span12Mux_h
    port map (
            O => \N__7182\,
            I => \N__7179\
        );

    \I__1283\ : Span12Mux_h
    port map (
            O => \N__7179\,
            I => \N__7176\
        );

    \I__1282\ : Odrv12
    port map (
            O => \N__7176\,
            I => mosi_output_c
        );

    \I__1281\ : InMux
    port map (
            O => \N__7173\,
            I => \N__7168\
        );

    \I__1280\ : InMux
    port map (
            O => \N__7172\,
            I => \N__7163\
        );

    \I__1279\ : InMux
    port map (
            O => \N__7171\,
            I => \N__7163\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__7168\,
            I => \switch_clk_2MHz_inst.aux_selection_2MHz_0\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__7163\,
            I => \switch_clk_2MHz_inst.aux_selection_2MHz_0\
        );

    \I__1276\ : InMux
    port map (
            O => \N__7158\,
            I => \N__7149\
        );

    \I__1275\ : InMux
    port map (
            O => \N__7157\,
            I => \N__7142\
        );

    \I__1274\ : InMux
    port map (
            O => \N__7156\,
            I => \N__7142\
        );

    \I__1273\ : InMux
    port map (
            O => \N__7155\,
            I => \N__7142\
        );

    \I__1272\ : InMux
    port map (
            O => \N__7154\,
            I => \N__7139\
        );

    \I__1271\ : InMux
    port map (
            O => \N__7153\,
            I => \N__7134\
        );

    \I__1270\ : InMux
    port map (
            O => \N__7152\,
            I => \N__7134\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__7149\,
            I => \switch_clk_2MHz_inst.N_91_li\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__7142\,
            I => \switch_clk_2MHz_inst.N_91_li\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__7139\,
            I => \switch_clk_2MHz_inst.N_91_li\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__7134\,
            I => \switch_clk_2MHz_inst.N_91_li\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__7125\,
            I => \switch_clk_2MHz_inst.SEL_0_RNI98MZ0Z31_cascade_\
        );

    \I__1264\ : CEMux
    port map (
            O => \N__7122\,
            I => \N__7119\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__7119\,
            I => \N_381_i\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__7116\,
            I => \switch_clk_2MHz_inst.counter_din_3_i_0_2_cascade_\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__7113\,
            I => \clk_out_RNI3LEM_cascade_\
        );

    \I__1260\ : InMux
    port map (
            O => \N__7110\,
            I => \N__7107\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__7107\,
            I => \switch_clk_2MHz_inst.G_31_0_o4_2\
        );

    \I__1258\ : InMux
    port map (
            O => \N__7104\,
            I => \N__7096\
        );

    \I__1257\ : InMux
    port map (
            O => \N__7103\,
            I => \N__7085\
        );

    \I__1256\ : InMux
    port map (
            O => \N__7102\,
            I => \N__7085\
        );

    \I__1255\ : InMux
    port map (
            O => \N__7101\,
            I => \N__7085\
        );

    \I__1254\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7085\
        );

    \I__1253\ : InMux
    port map (
            O => \N__7099\,
            I => \N__7085\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__7096\,
            I => \switch_clk_2MHz_inst.counter_dinZ0Z_0\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__7085\,
            I => \switch_clk_2MHz_inst.counter_dinZ0Z_0\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__7080\,
            I => \N__7074\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__7079\,
            I => \N__7071\
        );

    \I__1248\ : InMux
    port map (
            O => \N__7078\,
            I => \N__7067\
        );

    \I__1247\ : InMux
    port map (
            O => \N__7077\,
            I => \N__7064\
        );

    \I__1246\ : InMux
    port map (
            O => \N__7074\,
            I => \N__7057\
        );

    \I__1245\ : InMux
    port map (
            O => \N__7071\,
            I => \N__7057\
        );

    \I__1244\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7057\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__7067\,
            I => \switch_clk_2MHz_inst.counter_dinZ1Z_1\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__7064\,
            I => \switch_clk_2MHz_inst.counter_dinZ1Z_1\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__7057\,
            I => \switch_clk_2MHz_inst.counter_dinZ1Z_1\
        );

    \I__1240\ : InMux
    port map (
            O => \N__7050\,
            I => \N__7043\
        );

    \I__1239\ : InMux
    port map (
            O => \N__7049\,
            I => \N__7040\
        );

    \I__1238\ : InMux
    port map (
            O => \N__7048\,
            I => \N__7033\
        );

    \I__1237\ : InMux
    port map (
            O => \N__7047\,
            I => \N__7033\
        );

    \I__1236\ : InMux
    port map (
            O => \N__7046\,
            I => \N__7033\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__7043\,
            I => \switch_clk_2MHz_inst.counter_dinZ0Z_2\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__7040\,
            I => \switch_clk_2MHz_inst.counter_dinZ0Z_2\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__7033\,
            I => \switch_clk_2MHz_inst.counter_dinZ0Z_2\
        );

    \I__1232\ : InMux
    port map (
            O => \N__7026\,
            I => \N__7023\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__7023\,
            I => \switch_clk_2MHz_inst.N_92_0\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__7020\,
            I => \switch_clk_2MHz_inst.N_92_0_cascade_\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__7017\,
            I => \N__7012\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__7016\,
            I => \N__7009\
        );

    \I__1227\ : InMux
    port map (
            O => \N__7015\,
            I => \N__7006\
        );

    \I__1226\ : InMux
    port map (
            O => \N__7012\,
            I => \N__7003\
        );

    \I__1225\ : InMux
    port map (
            O => \N__7009\,
            I => \N__7000\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__7006\,
            I => \switch_clk_2MHz_inst.counter_dinZ0Z_3\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__7003\,
            I => \switch_clk_2MHz_inst.counter_dinZ0Z_3\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__7000\,
            I => \switch_clk_2MHz_inst.counter_dinZ0Z_3\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__6993\,
            I => \switch_clk_2MHz_inst.SEL_0_RNIC97QZ0_cascade_\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6990\,
            I => \N__6987\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6987\,
            I => \N__6984\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__6984\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_29\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6981\,
            I => \N__6978\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__6978\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_30\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6975\,
            I => \N__6972\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6972\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_83\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6969\,
            I => \N__6966\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6966\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_84\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6963\,
            I => \N__6960\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6960\,
            I => \N__6957\
        );

    \I__1209\ : Odrv4
    port map (
            O => \N__6957\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_41\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6954\,
            I => \N__6951\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6951\,
            I => \N__6948\
        );

    \I__1206\ : Odrv4
    port map (
            O => \N__6948\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_87\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__6945\,
            I => \N__6936\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6944\,
            I => \N__6913\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6943\,
            I => \N__6913\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6942\,
            I => \N__6913\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6941\,
            I => \N__6908\
        );

    \I__1200\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6908\
        );

    \I__1199\ : InMux
    port map (
            O => \N__6939\,
            I => \N__6905\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6936\,
            I => \N__6900\
        );

    \I__1197\ : InMux
    port map (
            O => \N__6935\,
            I => \N__6900\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6934\,
            I => \N__6893\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6933\,
            I => \N__6893\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6932\,
            I => \N__6893\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6931\,
            I => \N__6884\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6930\,
            I => \N__6884\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6929\,
            I => \N__6884\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6928\,
            I => \N__6884\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6927\,
            I => \N__6875\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6926\,
            I => \N__6866\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6866\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6924\,
            I => \N__6866\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6923\,
            I => \N__6866\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6922\,
            I => \N__6859\
        );

    \I__1183\ : InMux
    port map (
            O => \N__6921\,
            I => \N__6859\
        );

    \I__1182\ : InMux
    port map (
            O => \N__6920\,
            I => \N__6859\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6913\,
            I => \N__6855\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6908\,
            I => \N__6850\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6905\,
            I => \N__6850\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6900\,
            I => \N__6843\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6893\,
            I => \N__6843\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__6884\,
            I => \N__6843\
        );

    \I__1175\ : InMux
    port map (
            O => \N__6883\,
            I => \N__6836\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6882\,
            I => \N__6836\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6836\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6880\,
            I => \N__6829\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6879\,
            I => \N__6829\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6878\,
            I => \N__6829\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6875\,
            I => \N__6822\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6866\,
            I => \N__6822\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__6859\,
            I => \N__6822\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6858\,
            I => \N__6815\
        );

    \I__1165\ : Span4Mux_h
    port map (
            O => \N__6855\,
            I => \N__6810\
        );

    \I__1164\ : Span4Mux_h
    port map (
            O => \N__6850\,
            I => \N__6810\
        );

    \I__1163\ : Span4Mux_h
    port map (
            O => \N__6843\,
            I => \N__6807\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__6836\,
            I => \N__6802\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__6829\,
            I => \N__6802\
        );

    \I__1160\ : Span4Mux_h
    port map (
            O => \N__6822\,
            I => \N__6799\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6821\,
            I => \N__6794\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6820\,
            I => \N__6794\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6819\,
            I => \N__6789\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6818\,
            I => \N__6789\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6815\,
            I => \switch_clk_2MHz_inst.current_state_1_repZ0Z2\
        );

    \I__1154\ : Odrv4
    port map (
            O => \N__6810\,
            I => \switch_clk_2MHz_inst.current_state_1_repZ0Z2\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__6807\,
            I => \switch_clk_2MHz_inst.current_state_1_repZ0Z2\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__6802\,
            I => \switch_clk_2MHz_inst.current_state_1_repZ0Z2\
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__6799\,
            I => \switch_clk_2MHz_inst.current_state_1_repZ0Z2\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6794\,
            I => \switch_clk_2MHz_inst.current_state_1_repZ0Z2\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6789\,
            I => \switch_clk_2MHz_inst.current_state_1_repZ0Z2\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6771\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__6771\,
            I => \N__6768\
        );

    \I__1146\ : Odrv12
    port map (
            O => \N__6768\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_39\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6765\,
            I => \N__6762\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6762\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_40\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__6759\,
            I => \N__6747\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__6758\,
            I => \N__6740\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6757\,
            I => \N__6730\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6756\,
            I => \N__6730\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6755\,
            I => \N__6719\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6754\,
            I => \N__6719\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6753\,
            I => \N__6712\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6752\,
            I => \N__6712\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6751\,
            I => \N__6712\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6750\,
            I => \N__6707\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6747\,
            I => \N__6707\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6746\,
            I => \N__6702\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6745\,
            I => \N__6702\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6744\,
            I => \N__6691\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6743\,
            I => \N__6691\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6740\,
            I => \N__6691\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6739\,
            I => \N__6691\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6738\,
            I => \N__6691\
        );

    \I__1125\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6686\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6686\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__6735\,
            I => \N__6681\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__6730\,
            I => \N__6678\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6729\,
            I => \N__6665\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6728\,
            I => \N__6665\
        );

    \I__1119\ : InMux
    port map (
            O => \N__6727\,
            I => \N__6665\
        );

    \I__1118\ : InMux
    port map (
            O => \N__6726\,
            I => \N__6665\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6725\,
            I => \N__6660\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6724\,
            I => \N__6660\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__6719\,
            I => \N__6651\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6712\,
            I => \N__6651\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__6707\,
            I => \N__6651\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6702\,
            I => \N__6651\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__6691\,
            I => \N__6646\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6686\,
            I => \N__6646\
        );

    \I__1109\ : InMux
    port map (
            O => \N__6685\,
            I => \N__6641\
        );

    \I__1108\ : InMux
    port map (
            O => \N__6684\,
            I => \N__6641\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6681\,
            I => \N__6636\
        );

    \I__1106\ : Span12Mux_v
    port map (
            O => \N__6678\,
            I => \N__6633\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6677\,
            I => \N__6628\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6676\,
            I => \N__6628\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6623\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6623\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__6665\,
            I => \N__6618\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6660\,
            I => \N__6618\
        );

    \I__1099\ : Span4Mux_v
    port map (
            O => \N__6651\,
            I => \N__6611\
        );

    \I__1098\ : Span4Mux_s2_h
    port map (
            O => \N__6646\,
            I => \N__6611\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__6641\,
            I => \N__6611\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6606\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6639\,
            I => \N__6606\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6636\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_1\
        );

    \I__1093\ : Odrv12
    port map (
            O => \N__6633\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_1\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__6628\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_1\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__6623\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_1\
        );

    \I__1090\ : Odrv4
    port map (
            O => \N__6618\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_1\
        );

    \I__1089\ : Odrv4
    port map (
            O => \N__6611\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_1\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__6606\,
            I => \switch_clk_2MHz_inst.current_stateZ0Z_1\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6591\,
            I => \N__6588\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__6588\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_85\
        );

    \I__1085\ : InMux
    port map (
            O => \N__6585\,
            I => \N__6582\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__6582\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_86\
        );

    \I__1083\ : CEMux
    port map (
            O => \N__6579\,
            I => \N__6534\
        );

    \I__1082\ : CEMux
    port map (
            O => \N__6578\,
            I => \N__6534\
        );

    \I__1081\ : CEMux
    port map (
            O => \N__6577\,
            I => \N__6534\
        );

    \I__1080\ : CEMux
    port map (
            O => \N__6576\,
            I => \N__6534\
        );

    \I__1079\ : CEMux
    port map (
            O => \N__6575\,
            I => \N__6534\
        );

    \I__1078\ : CEMux
    port map (
            O => \N__6574\,
            I => \N__6534\
        );

    \I__1077\ : CEMux
    port map (
            O => \N__6573\,
            I => \N__6534\
        );

    \I__1076\ : CEMux
    port map (
            O => \N__6572\,
            I => \N__6534\
        );

    \I__1075\ : CEMux
    port map (
            O => \N__6571\,
            I => \N__6534\
        );

    \I__1074\ : CEMux
    port map (
            O => \N__6570\,
            I => \N__6534\
        );

    \I__1073\ : CEMux
    port map (
            O => \N__6569\,
            I => \N__6534\
        );

    \I__1072\ : CEMux
    port map (
            O => \N__6568\,
            I => \N__6534\
        );

    \I__1071\ : CEMux
    port map (
            O => \N__6567\,
            I => \N__6534\
        );

    \I__1070\ : CEMux
    port map (
            O => \N__6566\,
            I => \N__6534\
        );

    \I__1069\ : CEMux
    port map (
            O => \N__6565\,
            I => \N__6534\
        );

    \I__1068\ : GlobalMux
    port map (
            O => \N__6534\,
            I => \N__6531\
        );

    \I__1067\ : gio2CtrlBuf
    port map (
            O => \N__6531\,
            I => \switch_clk_2MHz_inst.N_259_g\
        );

    \I__1066\ : InMux
    port map (
            O => \N__6528\,
            I => \N__6525\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__6525\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_24\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6522\,
            I => \N__6519\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__6519\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_28\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__6516\,
            I => \N__6513\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6513\,
            I => \N__6510\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6510\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_57\
        );

    \I__1059\ : InMux
    port map (
            O => \N__6507\,
            I => \N__6504\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__6504\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_23\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6501\,
            I => \N__6498\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6498\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_27\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6495\,
            I => \N__6492\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__6492\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_25\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6489\,
            I => \N__6486\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6486\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_26\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6483\,
            I => \N__6480\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__6480\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_59\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6477\,
            I => \N__6474\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__6474\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_60\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6471\,
            I => \N__6468\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6468\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_61\
        );

    \I__1045\ : CascadeMux
    port map (
            O => \N__6465\,
            I => \switch_clk_1MHz_inst.current_state_cnv_0_1_cascade_\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6462\,
            I => \N__6458\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6461\,
            I => \N__6454\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6458\,
            I => \N__6451\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6457\,
            I => \N__6448\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6454\,
            I => \switch_clk_1MHz_inst.counter_dinZ1Z_1\
        );

    \I__1039\ : Odrv4
    port map (
            O => \N__6451\,
            I => \switch_clk_1MHz_inst.counter_dinZ1Z_1\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__6448\,
            I => \switch_clk_1MHz_inst.counter_dinZ1Z_1\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__6441\,
            I => \N__6437\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6440\,
            I => \N__6433\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6437\,
            I => \N__6427\
        );

    \I__1034\ : InMux
    port map (
            O => \N__6436\,
            I => \N__6427\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6433\,
            I => \N__6424\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6432\,
            I => \N__6421\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6427\,
            I => \switch_clk_1MHz_inst.counter_dinZ0Z_0\
        );

    \I__1030\ : Odrv4
    port map (
            O => \N__6424\,
            I => \switch_clk_1MHz_inst.counter_dinZ0Z_0\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6421\,
            I => \switch_clk_1MHz_inst.counter_dinZ0Z_0\
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__6414\,
            I => \switch_clk_1MHz_inst.current_state_RNO_8Z0Z_0_cascade_\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6411\,
            I => \N__6408\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__6408\,
            I => \switch_clk_1MHz_inst.current_state_RNO_2Z0Z_0\
        );

    \I__1025\ : CascadeMux
    port map (
            O => \N__6405\,
            I => \N__6402\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6402\,
            I => \N__6395\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6401\,
            I => \N__6395\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6400\,
            I => \N__6392\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__6395\,
            I => \switch_clk_1MHz_inst.N_88_0\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__6392\,
            I => \switch_clk_1MHz_inst.N_88_0\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6387\,
            I => \N__6383\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6386\,
            I => \N__6378\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__6383\,
            I => \N__6375\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6382\,
            I => \N__6370\
        );

    \I__1015\ : InMux
    port map (
            O => \N__6381\,
            I => \N__6370\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__6378\,
            I => \switch_clk_1MHz_inst.counter_dinZ0Z_2\
        );

    \I__1013\ : Odrv4
    port map (
            O => \N__6375\,
            I => \switch_clk_1MHz_inst.counter_dinZ0Z_2\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6370\,
            I => \switch_clk_1MHz_inst.counter_dinZ0Z_2\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6363\,
            I => \N__6360\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__6360\,
            I => \switch_clk_2MHz_inst.N_8_0\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6348\
        );

    \I__1008\ : InMux
    port map (
            O => \N__6356\,
            I => \N__6348\
        );

    \I__1007\ : InMux
    port map (
            O => \N__6355\,
            I => \N__6348\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6348\,
            I => \N__6341\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6347\,
            I => \N__6332\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6346\,
            I => \N__6332\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6345\,
            I => \N__6332\
        );

    \I__1002\ : InMux
    port map (
            O => \N__6344\,
            I => \N__6332\
        );

    \I__1001\ : Odrv4
    port map (
            O => \N__6341\,
            I => \switch_clk_1MHz_inst.current_state_d_i_2\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__6332\,
            I => \switch_clk_1MHz_inst.current_state_d_i_2\
        );

    \I__999\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6311\
        );

    \I__998\ : InMux
    port map (
            O => \N__6326\,
            I => \N__6311\
        );

    \I__997\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6311\
        );

    \I__996\ : InMux
    port map (
            O => \N__6324\,
            I => \N__6311\
        );

    \I__995\ : InMux
    port map (
            O => \N__6323\,
            I => \N__6302\
        );

    \I__994\ : InMux
    port map (
            O => \N__6322\,
            I => \N__6302\
        );

    \I__993\ : InMux
    port map (
            O => \N__6321\,
            I => \N__6302\
        );

    \I__992\ : InMux
    port map (
            O => \N__6320\,
            I => \N__6302\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__6311\,
            I => \switch_clk_1MHz_inst.N_116_1_i\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__6302\,
            I => \switch_clk_1MHz_inst.N_116_1_i\
        );

    \I__989\ : InMux
    port map (
            O => \N__6297\,
            I => \N__6294\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__6294\,
            I => \N__6291\
        );

    \I__987\ : Span12Mux_s10_v
    port map (
            O => \N__6291\,
            I => \N__6288\
        );

    \I__986\ : Odrv12
    port map (
            O => \N__6288\,
            I => \config_register_latched_dec_inst.DYNCNF_0\
        );

    \I__985\ : InMux
    port map (
            O => \N__6285\,
            I => \N__6279\
        );

    \I__984\ : InMux
    port map (
            O => \N__6284\,
            I => \N__6279\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__6279\,
            I => \config_register_latched_dec_inst.DYNCNF_1Z0Z_0\
        );

    \I__982\ : CascadeMux
    port map (
            O => \N__6276\,
            I => \counter_RNISR1F_2_cascade_\
        );

    \I__981\ : IoInMux
    port map (
            O => \N__6273\,
            I => \N__6270\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__6270\,
            I => \N__6267\
        );

    \I__979\ : Span12Mux_s2_v
    port map (
            O => \N__6267\,
            I => \N__6264\
        );

    \I__978\ : Span12Mux_h
    port map (
            O => \N__6264\,
            I => \N__6261\
        );

    \I__977\ : Odrv12
    port map (
            O => \N__6261\,
            I => \switch_clk_1MHz_inst.current_state_RNITOE91_0Z0Z_1\
        );

    \I__976\ : InMux
    port map (
            O => \N__6258\,
            I => \N__6253\
        );

    \I__975\ : InMux
    port map (
            O => \N__6257\,
            I => \N__6250\
        );

    \I__974\ : InMux
    port map (
            O => \N__6256\,
            I => \N__6247\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__6253\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_3\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__6250\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_3\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__6247\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_3\
        );

    \I__970\ : InMux
    port map (
            O => \N__6240\,
            I => \N__6223\
        );

    \I__969\ : InMux
    port map (
            O => \N__6239\,
            I => \N__6223\
        );

    \I__968\ : InMux
    port map (
            O => \N__6238\,
            I => \N__6223\
        );

    \I__967\ : InMux
    port map (
            O => \N__6237\,
            I => \N__6223\
        );

    \I__966\ : InMux
    port map (
            O => \N__6236\,
            I => \N__6220\
        );

    \I__965\ : InMux
    port map (
            O => \N__6235\,
            I => \N__6213\
        );

    \I__964\ : InMux
    port map (
            O => \N__6234\,
            I => \N__6213\
        );

    \I__963\ : InMux
    port map (
            O => \N__6233\,
            I => \N__6213\
        );

    \I__962\ : CascadeMux
    port map (
            O => \N__6232\,
            I => \N__6210\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__6223\,
            I => \N__6206\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__6220\,
            I => \N__6201\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__6213\,
            I => \N__6201\
        );

    \I__958\ : InMux
    port map (
            O => \N__6210\,
            I => \N__6198\
        );

    \I__957\ : InMux
    port map (
            O => \N__6209\,
            I => \N__6195\
        );

    \I__956\ : Span4Mux_v
    port map (
            O => \N__6206\,
            I => \N__6190\
        );

    \I__955\ : Span4Mux_v
    port map (
            O => \N__6201\,
            I => \N__6190\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__6198\,
            I => \switch_clk_2MHz_inst.current_state_fastZ0Z_1\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__6195\,
            I => \switch_clk_2MHz_inst.current_state_fastZ0Z_1\
        );

    \I__952\ : Odrv4
    port map (
            O => \N__6190\,
            I => \switch_clk_2MHz_inst.current_state_fastZ0Z_1\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__6183\,
            I => \switch_clk_2MHz_inst.counter_statlde_0_cascade_\
        );

    \I__950\ : CEMux
    port map (
            O => \N__6180\,
            I => \N__6177\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__6177\,
            I => \N__6174\
        );

    \I__948\ : Odrv4
    port map (
            O => \N__6174\,
            I => \switch_clk_2MHz_inst.current_state_fast_RNI9DAU1Z0Z_1\
        );

    \I__947\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6167\
        );

    \I__946\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6164\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__6167\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_1\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__6164\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_1\
        );

    \I__943\ : InMux
    port map (
            O => \N__6159\,
            I => \N__6154\
        );

    \I__942\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6149\
        );

    \I__941\ : InMux
    port map (
            O => \N__6157\,
            I => \N__6149\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__6154\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_6\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__6149\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_6\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__6144\,
            I => \N__6140\
        );

    \I__937\ : InMux
    port map (
            O => \N__6143\,
            I => \N__6136\
        );

    \I__936\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6133\
        );

    \I__935\ : InMux
    port map (
            O => \N__6139\,
            I => \N__6130\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__6136\,
            I => \N__6125\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__6133\,
            I => \N__6125\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__6130\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_5\
        );

    \I__931\ : Odrv4
    port map (
            O => \N__6125\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_5\
        );

    \I__930\ : InMux
    port map (
            O => \N__6120\,
            I => \N__6113\
        );

    \I__929\ : InMux
    port map (
            O => \N__6119\,
            I => \N__6113\
        );

    \I__928\ : InMux
    port map (
            O => \N__6118\,
            I => \N__6110\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__6113\,
            I => \N__6107\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__6110\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_4\
        );

    \I__925\ : Odrv4
    port map (
            O => \N__6107\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_4\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__6102\,
            I => \switch_clk_2MHz_inst.G_31_0_a4_1_1_cascade_\
        );

    \I__923\ : InMux
    port map (
            O => \N__6099\,
            I => \N__6096\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__6096\,
            I => \switch_clk_2MHz_inst.G_31_0_a4_1_5\
        );

    \I__921\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6090\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__6090\,
            I => \switch_clk_2MHz_inst.N_9_1\
        );

    \I__919\ : CascadeMux
    port map (
            O => \N__6087\,
            I => \switch_clk_2MHz_inst.G_31_0_a4_1_6_cascade_\
        );

    \I__918\ : InMux
    port map (
            O => \N__6084\,
            I => \N__6080\
        );

    \I__917\ : InMux
    port map (
            O => \N__6083\,
            I => \N__6077\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__6080\,
            I => \N__6074\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__6077\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_2\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__6074\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_2\
        );

    \I__913\ : InMux
    port map (
            O => \N__6069\,
            I => \N__6065\
        );

    \I__912\ : InMux
    port map (
            O => \N__6068\,
            I => \N__6062\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__6065\,
            I => \N__6059\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__6062\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_1\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__6059\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_1\
        );

    \I__908\ : CascadeMux
    port map (
            O => \N__6054\,
            I => \N__6051\
        );

    \I__907\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6046\
        );

    \I__906\ : InMux
    port map (
            O => \N__6050\,
            I => \N__6043\
        );

    \I__905\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6040\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__6046\,
            I => \N__6037\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__6043\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_5\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__6040\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_5\
        );

    \I__901\ : Odrv4
    port map (
            O => \N__6037\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_5\
        );

    \I__900\ : InMux
    port map (
            O => \N__6030\,
            I => \N__6026\
        );

    \I__899\ : InMux
    port map (
            O => \N__6029\,
            I => \N__6023\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__6026\,
            I => \N__6020\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__6023\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_0\
        );

    \I__896\ : Odrv4
    port map (
            O => \N__6020\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_0\
        );

    \I__895\ : InMux
    port map (
            O => \N__6015\,
            I => \N__6012\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__6012\,
            I => \N__6009\
        );

    \I__893\ : Span4Mux_v
    port map (
            O => \N__6009\,
            I => \N__6006\
        );

    \I__892\ : Odrv4
    port map (
            O => \N__6006\,
            I => \switch_clk_1MHz_inst.current_state_RNO_3Z0Z_0\
        );

    \I__891\ : InMux
    port map (
            O => \N__6003\,
            I => \N__5998\
        );

    \I__890\ : InMux
    port map (
            O => \N__6002\,
            I => \N__5995\
        );

    \I__889\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5992\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5998\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_4\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5995\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_4\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__5992\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_4\
        );

    \I__885\ : InMux
    port map (
            O => \N__5985\,
            I => \N__5981\
        );

    \I__884\ : InMux
    port map (
            O => \N__5984\,
            I => \N__5978\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__5981\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_1\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__5978\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_1\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__5973\,
            I => \N__5968\
        );

    \I__880\ : InMux
    port map (
            O => \N__5972\,
            I => \N__5965\
        );

    \I__879\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5962\
        );

    \I__878\ : InMux
    port map (
            O => \N__5968\,
            I => \N__5959\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5965\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_5\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5962\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_5\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5959\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_5\
        );

    \I__874\ : InMux
    port map (
            O => \N__5952\,
            I => \N__5949\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5949\,
            I => \switch_clk_1MHz_inst.current_state_ns_0_a3_1_5_0\
        );

    \I__872\ : CascadeMux
    port map (
            O => \N__5946\,
            I => \N__5943\
        );

    \I__871\ : InMux
    port map (
            O => \N__5943\,
            I => \N__5940\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5940\,
            I => \N__5937\
        );

    \I__869\ : Span4Mux_h
    port map (
            O => \N__5937\,
            I => \N__5934\
        );

    \I__868\ : Odrv4
    port map (
            O => \N__5934\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_15\
        );

    \I__867\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5928\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5928\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_47\
        );

    \I__865\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5922\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5922\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_48\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__5919\,
            I => \N__5916\
        );

    \I__862\ : InMux
    port map (
            O => \N__5916\,
            I => \N__5913\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5913\,
            I => \N__5910\
        );

    \I__860\ : Odrv4
    port map (
            O => \N__5910\,
            I => \switch_clk_2MHz_inst.flag_input_regZ0\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__5907\,
            I => \switch_clk_2MHz_inst.N_114_0_cascade_\
        );

    \I__858\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5897\
        );

    \I__857\ : InMux
    port map (
            O => \N__5903\,
            I => \N__5897\
        );

    \I__856\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5894\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__5897\,
            I => \N__5867\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__5894\,
            I => \N__5867\
        );

    \I__853\ : InMux
    port map (
            O => \N__5893\,
            I => \N__5856\
        );

    \I__852\ : InMux
    port map (
            O => \N__5892\,
            I => \N__5856\
        );

    \I__851\ : InMux
    port map (
            O => \N__5891\,
            I => \N__5856\
        );

    \I__850\ : InMux
    port map (
            O => \N__5890\,
            I => \N__5856\
        );

    \I__849\ : InMux
    port map (
            O => \N__5889\,
            I => \N__5856\
        );

    \I__848\ : InMux
    port map (
            O => \N__5888\,
            I => \N__5843\
        );

    \I__847\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5843\
        );

    \I__846\ : InMux
    port map (
            O => \N__5886\,
            I => \N__5843\
        );

    \I__845\ : InMux
    port map (
            O => \N__5885\,
            I => \N__5843\
        );

    \I__844\ : InMux
    port map (
            O => \N__5884\,
            I => \N__5843\
        );

    \I__843\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5843\
        );

    \I__842\ : InMux
    port map (
            O => \N__5882\,
            I => \N__5838\
        );

    \I__841\ : InMux
    port map (
            O => \N__5881\,
            I => \N__5838\
        );

    \I__840\ : InMux
    port map (
            O => \N__5880\,
            I => \N__5833\
        );

    \I__839\ : InMux
    port map (
            O => \N__5879\,
            I => \N__5833\
        );

    \I__838\ : InMux
    port map (
            O => \N__5878\,
            I => \N__5828\
        );

    \I__837\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5823\
        );

    \I__836\ : InMux
    port map (
            O => \N__5876\,
            I => \N__5823\
        );

    \I__835\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5820\
        );

    \I__834\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5813\
        );

    \I__833\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5813\
        );

    \I__832\ : InMux
    port map (
            O => \N__5872\,
            I => \N__5813\
        );

    \I__831\ : Span4Mux_v
    port map (
            O => \N__5867\,
            I => \N__5806\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5856\,
            I => \N__5806\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__5843\,
            I => \N__5806\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5838\,
            I => \N__5801\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__5833\,
            I => \N__5801\
        );

    \I__826\ : InMux
    port map (
            O => \N__5832\,
            I => \N__5798\
        );

    \I__825\ : InMux
    port map (
            O => \N__5831\,
            I => \N__5789\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5828\,
            I => \N__5784\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__5823\,
            I => \N__5784\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5820\,
            I => \N__5781\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5813\,
            I => \N__5778\
        );

    \I__820\ : Span4Mux_v
    port map (
            O => \N__5806\,
            I => \N__5774\
        );

    \I__819\ : Span4Mux_h
    port map (
            O => \N__5801\,
            I => \N__5771\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5798\,
            I => \N__5768\
        );

    \I__817\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5755\
        );

    \I__816\ : InMux
    port map (
            O => \N__5796\,
            I => \N__5755\
        );

    \I__815\ : InMux
    port map (
            O => \N__5795\,
            I => \N__5755\
        );

    \I__814\ : InMux
    port map (
            O => \N__5794\,
            I => \N__5755\
        );

    \I__813\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5755\
        );

    \I__812\ : InMux
    port map (
            O => \N__5792\,
            I => \N__5755\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__5789\,
            I => \N__5746\
        );

    \I__810\ : Span4Mux_v
    port map (
            O => \N__5784\,
            I => \N__5746\
        );

    \I__809\ : Span4Mux_s3_h
    port map (
            O => \N__5781\,
            I => \N__5746\
        );

    \I__808\ : Span4Mux_s3_h
    port map (
            O => \N__5778\,
            I => \N__5746\
        );

    \I__807\ : InMux
    port map (
            O => \N__5777\,
            I => \N__5743\
        );

    \I__806\ : Odrv4
    port map (
            O => \N__5774\,
            I => \switch_clk_2MHz_inst.current_state_1_repZ0Z1\
        );

    \I__805\ : Odrv4
    port map (
            O => \N__5771\,
            I => \switch_clk_2MHz_inst.current_state_1_repZ0Z1\
        );

    \I__804\ : Odrv4
    port map (
            O => \N__5768\,
            I => \switch_clk_2MHz_inst.current_state_1_repZ0Z1\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5755\,
            I => \switch_clk_2MHz_inst.current_state_1_repZ0Z1\
        );

    \I__802\ : Odrv4
    port map (
            O => \N__5746\,
            I => \switch_clk_2MHz_inst.current_state_1_repZ0Z1\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5743\,
            I => \switch_clk_2MHz_inst.current_state_1_repZ0Z1\
        );

    \I__800\ : InMux
    port map (
            O => \N__5730\,
            I => \N__5717\
        );

    \I__799\ : InMux
    port map (
            O => \N__5729\,
            I => \N__5717\
        );

    \I__798\ : InMux
    port map (
            O => \N__5728\,
            I => \N__5717\
        );

    \I__797\ : InMux
    port map (
            O => \N__5727\,
            I => \N__5708\
        );

    \I__796\ : InMux
    port map (
            O => \N__5726\,
            I => \N__5708\
        );

    \I__795\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5708\
        );

    \I__794\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5708\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__5717\,
            I => \switch_clk_2MHz_inst.current_state_d_i_2\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5708\,
            I => \switch_clk_2MHz_inst.current_state_d_i_2\
        );

    \I__791\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5700\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5700\,
            I => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_58\
        );

    \I__789\ : IoInMux
    port map (
            O => \N__5697\,
            I => \N__5694\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__5694\,
            I => \N__5691\
        );

    \I__787\ : Span4Mux_s0_v
    port map (
            O => \N__5691\,
            I => \N__5688\
        );

    \I__786\ : Span4Mux_v
    port map (
            O => \N__5688\,
            I => \N__5685\
        );

    \I__785\ : Odrv4
    port map (
            O => \N__5685\,
            I => \DYNCNF_i_0\
        );

    \I__784\ : InMux
    port map (
            O => \N__5682\,
            I => \N__5679\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5679\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_82\
        );

    \I__782\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5673\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5673\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_61\
        );

    \I__780\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5667\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5667\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_46\
        );

    \I__778\ : InMux
    port map (
            O => \N__5664\,
            I => \N__5661\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5661\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_59\
        );

    \I__776\ : InMux
    port map (
            O => \N__5658\,
            I => \N__5655\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5655\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_60\
        );

    \I__774\ : InMux
    port map (
            O => \N__5652\,
            I => \switch_clk_1MHz_inst.counter_idle_cry_5\
        );

    \I__773\ : InMux
    port map (
            O => \N__5649\,
            I => \switch_clk_1MHz_inst.counter_idle_cry_6\
        );

    \I__772\ : InMux
    port map (
            O => \N__5646\,
            I => \N__5643\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5643\,
            I => \switch_clk_1MHz_inst.N_116_1\
        );

    \I__770\ : CascadeMux
    port map (
            O => \N__5640\,
            I => \switch_clk_1MHz_inst.G_31_1_cascade_\
        );

    \I__769\ : CEMux
    port map (
            O => \N__5637\,
            I => \N__5634\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5634\,
            I => \switch_clk_1MHz_inst.counter_idle_RNIOJRU1Z0Z_7\
        );

    \I__767\ : InMux
    port map (
            O => \N__5631\,
            I => \N__5626\
        );

    \I__766\ : InMux
    port map (
            O => \N__5630\,
            I => \N__5621\
        );

    \I__765\ : InMux
    port map (
            O => \N__5629\,
            I => \N__5621\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5626\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_3\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__5621\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_3\
        );

    \I__762\ : InMux
    port map (
            O => \N__5616\,
            I => \N__5611\
        );

    \I__761\ : InMux
    port map (
            O => \N__5615\,
            I => \N__5606\
        );

    \I__760\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5606\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5611\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_4\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5606\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_4\
        );

    \I__757\ : InMux
    port map (
            O => \N__5601\,
            I => \N__5594\
        );

    \I__756\ : InMux
    port map (
            O => \N__5600\,
            I => \N__5594\
        );

    \I__755\ : InMux
    port map (
            O => \N__5599\,
            I => \N__5591\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5594\,
            I => \N__5588\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__5591\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_7\
        );

    \I__752\ : Odrv4
    port map (
            O => \N__5588\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_7\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__5583\,
            I => \N__5579\
        );

    \I__750\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5573\
        );

    \I__749\ : InMux
    port map (
            O => \N__5579\,
            I => \N__5573\
        );

    \I__748\ : InMux
    port map (
            O => \N__5578\,
            I => \N__5570\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__5573\,
            I => \N__5567\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__5570\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_6\
        );

    \I__745\ : Odrv4
    port map (
            O => \N__5567\,
            I => \switch_clk_1MHz_inst.counter_idleZ0Z_6\
        );

    \I__744\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5559\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__5559\,
            I => \switch_clk_1MHz_inst.current_state_RNO_5Z0Z_0\
        );

    \I__742\ : CascadeMux
    port map (
            O => \N__5556\,
            I => \switch_clk_1MHz_inst.current_state_RNO_4Z0Z_0_cascade_\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__5553\,
            I => \switch_clk_1MHz_inst.N_116_cascade_\
        );

    \I__740\ : InMux
    port map (
            O => \N__5550\,
            I => \N__5547\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__5547\,
            I => \N__5544\
        );

    \I__738\ : Odrv4
    port map (
            O => \N__5544\,
            I => \switch_clk_1MHz_inst.current_state_RNO_1Z0Z_0\
        );

    \I__737\ : InMux
    port map (
            O => \N__5541\,
            I => \switch_clk_1MHz_inst.counter_stat_cry_3\
        );

    \I__736\ : InMux
    port map (
            O => \N__5538\,
            I => \switch_clk_1MHz_inst.counter_stat_cry_4\
        );

    \I__735\ : InMux
    port map (
            O => \N__5535\,
            I => \switch_clk_1MHz_inst.counter_stat_cry_5\
        );

    \I__734\ : CascadeMux
    port map (
            O => \N__5532\,
            I => \N__5527\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__5531\,
            I => \N__5524\
        );

    \I__732\ : InMux
    port map (
            O => \N__5530\,
            I => \N__5521\
        );

    \I__731\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5518\
        );

    \I__730\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5515\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__5521\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_6\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__5518\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_6\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__5515\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_6\
        );

    \I__726\ : CEMux
    port map (
            O => \N__5508\,
            I => \N__5505\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5505\,
            I => \N__5502\
        );

    \I__724\ : Span4Mux_v
    port map (
            O => \N__5502\,
            I => \N__5499\
        );

    \I__723\ : Span4Mux_s3_h
    port map (
            O => \N__5499\,
            I => \N__5496\
        );

    \I__722\ : Odrv4
    port map (
            O => \N__5496\,
            I => \switch_clk_1MHz_inst.current_state_RNIFA8B2Z0Z_1\
        );

    \I__721\ : InMux
    port map (
            O => \N__5493\,
            I => \bfn_4_23_0_\
        );

    \I__720\ : InMux
    port map (
            O => \N__5490\,
            I => \switch_clk_1MHz_inst.counter_idle_cry_0\
        );

    \I__719\ : InMux
    port map (
            O => \N__5487\,
            I => \switch_clk_1MHz_inst.counter_idle_cry_1\
        );

    \I__718\ : InMux
    port map (
            O => \N__5484\,
            I => \switch_clk_1MHz_inst.counter_idle_cry_2\
        );

    \I__717\ : InMux
    port map (
            O => \N__5481\,
            I => \switch_clk_1MHz_inst.counter_idle_cry_3\
        );

    \I__716\ : InMux
    port map (
            O => \N__5478\,
            I => \switch_clk_1MHz_inst.counter_idle_cry_4\
        );

    \I__715\ : InMux
    port map (
            O => \N__5475\,
            I => \N__5470\
        );

    \I__714\ : InMux
    port map (
            O => \N__5474\,
            I => \N__5467\
        );

    \I__713\ : InMux
    port map (
            O => \N__5473\,
            I => \N__5464\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__5470\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_4\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__5467\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_4\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5464\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_4\
        );

    \I__709\ : InMux
    port map (
            O => \N__5457\,
            I => \N__5452\
        );

    \I__708\ : InMux
    port map (
            O => \N__5456\,
            I => \N__5449\
        );

    \I__707\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5446\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5452\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_3\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__5449\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_3\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5446\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_3\
        );

    \I__703\ : InMux
    port map (
            O => \N__5439\,
            I => \N__5436\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5436\,
            I => \switch_clk_2MHz_inst.G_31_0_a4_0_4\
        );

    \I__701\ : CascadeMux
    port map (
            O => \N__5433\,
            I => \switch_clk_2MHz_inst.G_31_0_a4_0_5_cascade_\
        );

    \I__700\ : CascadeMux
    port map (
            O => \N__5430\,
            I => \switch_clk_1MHz_inst.current_state_ns_0_a3_1_4_0_cascade_\
        );

    \I__699\ : InMux
    port map (
            O => \N__5427\,
            I => \N__5415\
        );

    \I__698\ : InMux
    port map (
            O => \N__5426\,
            I => \N__5415\
        );

    \I__697\ : InMux
    port map (
            O => \N__5425\,
            I => \N__5415\
        );

    \I__696\ : InMux
    port map (
            O => \N__5424\,
            I => \N__5408\
        );

    \I__695\ : InMux
    port map (
            O => \N__5423\,
            I => \N__5408\
        );

    \I__694\ : InMux
    port map (
            O => \N__5422\,
            I => \N__5408\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__5415\,
            I => \switch_clk_2MHz_inst.N_117_1_i\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5408\,
            I => \switch_clk_2MHz_inst.N_117_1_i\
        );

    \I__691\ : InMux
    port map (
            O => \N__5403\,
            I => \N__5399\
        );

    \I__690\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5396\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5399\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_0\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__5396\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_0\
        );

    \I__687\ : InMux
    port map (
            O => \N__5391\,
            I => \bfn_4_22_0_\
        );

    \I__686\ : InMux
    port map (
            O => \N__5388\,
            I => \switch_clk_1MHz_inst.counter_stat_cry_0\
        );

    \I__685\ : InMux
    port map (
            O => \N__5385\,
            I => \N__5381\
        );

    \I__684\ : InMux
    port map (
            O => \N__5384\,
            I => \N__5378\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__5381\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_2\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5378\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_2\
        );

    \I__681\ : InMux
    port map (
            O => \N__5373\,
            I => \switch_clk_1MHz_inst.counter_stat_cry_1\
        );

    \I__680\ : InMux
    port map (
            O => \N__5370\,
            I => \N__5365\
        );

    \I__679\ : InMux
    port map (
            O => \N__5369\,
            I => \N__5362\
        );

    \I__678\ : InMux
    port map (
            O => \N__5368\,
            I => \N__5359\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__5365\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_3\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__5362\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_3\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__5359\,
            I => \switch_clk_1MHz_inst.counter_statZ0Z_3\
        );

    \I__674\ : InMux
    port map (
            O => \N__5352\,
            I => \switch_clk_1MHz_inst.counter_stat_cry_2\
        );

    \I__673\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5346\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__5346\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_5\
        );

    \I__671\ : CascadeMux
    port map (
            O => \N__5343\,
            I => \N__5340\
        );

    \I__670\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5337\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5337\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_6\
        );

    \I__668\ : InMux
    port map (
            O => \N__5334\,
            I => \N__5330\
        );

    \I__667\ : InMux
    port map (
            O => \N__5333\,
            I => \N__5327\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__5330\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_0\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__5327\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_0\
        );

    \I__664\ : InMux
    port map (
            O => \N__5322\,
            I => \bfn_4_20_0_\
        );

    \I__663\ : InMux
    port map (
            O => \N__5319\,
            I => \switch_clk_2MHz_inst.counter_stat_cry_0\
        );

    \I__662\ : CascadeMux
    port map (
            O => \N__5316\,
            I => \N__5313\
        );

    \I__661\ : InMux
    port map (
            O => \N__5313\,
            I => \N__5309\
        );

    \I__660\ : InMux
    port map (
            O => \N__5312\,
            I => \N__5306\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__5309\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_2\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__5306\,
            I => \switch_clk_2MHz_inst.counter_statZ0Z_2\
        );

    \I__657\ : InMux
    port map (
            O => \N__5301\,
            I => \switch_clk_2MHz_inst.counter_stat_cry_1\
        );

    \I__656\ : InMux
    port map (
            O => \N__5298\,
            I => \switch_clk_2MHz_inst.counter_stat_cry_2\
        );

    \I__655\ : InMux
    port map (
            O => \N__5295\,
            I => \switch_clk_2MHz_inst.counter_stat_cry_3\
        );

    \I__654\ : InMux
    port map (
            O => \N__5292\,
            I => \switch_clk_2MHz_inst.counter_stat_cry_4\
        );

    \I__653\ : InMux
    port map (
            O => \N__5289\,
            I => \switch_clk_2MHz_inst.counter_stat_cry_5\
        );

    \I__652\ : InMux
    port map (
            O => \N__5286\,
            I => \N__5282\
        );

    \I__651\ : InMux
    port map (
            O => \N__5285\,
            I => \N__5279\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__5282\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_0\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__5279\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_0\
        );

    \I__648\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5270\
        );

    \I__647\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5267\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__5270\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_1\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__5267\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_1\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__5262\,
            I => \N__5257\
        );

    \I__643\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5254\
        );

    \I__642\ : InMux
    port map (
            O => \N__5260\,
            I => \N__5251\
        );

    \I__641\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5248\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__5254\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_2\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__5251\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_2\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__5248\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_2\
        );

    \I__637\ : CascadeMux
    port map (
            O => \N__5241\,
            I => \N__5236\
        );

    \I__636\ : InMux
    port map (
            O => \N__5240\,
            I => \N__5233\
        );

    \I__635\ : InMux
    port map (
            O => \N__5239\,
            I => \N__5230\
        );

    \I__634\ : InMux
    port map (
            O => \N__5236\,
            I => \N__5227\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__5233\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_5\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__5230\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_5\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__5227\,
            I => \switch_clk_2MHz_inst.counter_idleZ0Z_5\
        );

    \I__630\ : InMux
    port map (
            O => \N__5220\,
            I => \N__5217\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__5217\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_49\
        );

    \I__628\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5211\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__5211\,
            I => \N__5208\
        );

    \I__626\ : Odrv4
    port map (
            O => \N__5208\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_45\
        );

    \I__625\ : InMux
    port map (
            O => \N__5205\,
            I => \N__5202\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__5202\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_7\
        );

    \I__623\ : InMux
    port map (
            O => \N__5199\,
            I => \N__5196\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__5196\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_24\
        );

    \I__621\ : InMux
    port map (
            O => \N__5193\,
            I => \N__5190\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__5190\,
            I => \N__5187\
        );

    \I__619\ : Odrv4
    port map (
            O => \N__5187\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_25\
        );

    \I__618\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5181\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__5181\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_3\
        );

    \I__616\ : InMux
    port map (
            O => \N__5178\,
            I => \N__5175\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__5175\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_0\
        );

    \I__614\ : InMux
    port map (
            O => \N__5172\,
            I => \N__5169\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__5169\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_1\
        );

    \I__612\ : InMux
    port map (
            O => \N__5166\,
            I => \N__5163\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__5163\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_2\
        );

    \I__610\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5157\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__5157\,
            I => \N__5154\
        );

    \I__608\ : Odrv4
    port map (
            O => \N__5154\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_69\
        );

    \I__607\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5148\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__5148\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_70\
        );

    \I__605\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5142\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__5142\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_71\
        );

    \I__603\ : InMux
    port map (
            O => \N__5139\,
            I => \N__5136\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__5136\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_22\
        );

    \I__601\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5130\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__5130\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_62\
        );

    \I__599\ : InMux
    port map (
            O => \N__5127\,
            I => \N__5124\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__5124\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_63\
        );

    \I__597\ : InMux
    port map (
            O => \N__5121\,
            I => \N__5118\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__5118\,
            I => \N__5115\
        );

    \I__595\ : Odrv4
    port map (
            O => \N__5115\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_58\
        );

    \I__594\ : InMux
    port map (
            O => \N__5112\,
            I => \N__5109\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__5109\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_23\
        );

    \I__592\ : InMux
    port map (
            O => \N__5106\,
            I => \N__5103\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__5103\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_4\
        );

    \I__590\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5097\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__5097\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_10\
        );

    \I__588\ : InMux
    port map (
            O => \N__5094\,
            I => \N__5091\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__5091\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_11\
        );

    \I__586\ : InMux
    port map (
            O => \N__5088\,
            I => \N__5085\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__5085\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_14\
        );

    \I__584\ : InMux
    port map (
            O => \N__5082\,
            I => \N__5079\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__5079\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_12\
        );

    \I__582\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5073\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__5073\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_13\
        );

    \I__580\ : CascadeMux
    port map (
            O => \N__5070\,
            I => \switch_clk_1MHz_inst.counter_statlde_0_cascade_\
        );

    \I__579\ : CEMux
    port map (
            O => \N__5067\,
            I => \N__5062\
        );

    \I__578\ : CEMux
    port map (
            O => \N__5066\,
            I => \N__5059\
        );

    \I__577\ : CEMux
    port map (
            O => \N__5065\,
            I => \N__5056\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__5062\,
            I => \switch_clk_1MHz_inst.current_state_RNITOE91Z0Z_1\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__5059\,
            I => \switch_clk_1MHz_inst.current_state_RNITOE91Z0Z_1\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__5056\,
            I => \switch_clk_1MHz_inst.current_state_RNITOE91Z0Z_1\
        );

    \I__573\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5046\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__5046\,
            I => \N__5043\
        );

    \I__571\ : Odrv4
    port map (
            O => \N__5043\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_72\
        );

    \I__570\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5037\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__5037\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_81\
        );

    \I__568\ : InMux
    port map (
            O => \N__5034\,
            I => \bfn_3_21_0_\
        );

    \I__567\ : InMux
    port map (
            O => \N__5031\,
            I => \switch_clk_2MHz_inst.counter_idle_cry_0\
        );

    \I__566\ : InMux
    port map (
            O => \N__5028\,
            I => \switch_clk_2MHz_inst.counter_idle_cry_1\
        );

    \I__565\ : InMux
    port map (
            O => \N__5025\,
            I => \switch_clk_2MHz_inst.counter_idle_cry_2\
        );

    \I__564\ : InMux
    port map (
            O => \N__5022\,
            I => \switch_clk_2MHz_inst.counter_idle_cry_3\
        );

    \I__563\ : InMux
    port map (
            O => \N__5019\,
            I => \switch_clk_2MHz_inst.counter_idle_cry_4\
        );

    \I__562\ : CEMux
    port map (
            O => \N__5016\,
            I => \N__5013\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__5013\,
            I => \N__5010\
        );

    \I__560\ : Span4Mux_h
    port map (
            O => \N__5010\,
            I => \N__5007\
        );

    \I__559\ : Odrv4
    port map (
            O => \N__5007\,
            I => \switch_clk_2MHz_inst.current_state_fast_RNIDHKD1Z0Z_1\
        );

    \I__558\ : InMux
    port map (
            O => \N__5004\,
            I => \N__5001\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__5001\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_8\
        );

    \I__556\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4995\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4995\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_9\
        );

    \I__554\ : InMux
    port map (
            O => \N__4992\,
            I => \N__4989\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__4989\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_33\
        );

    \I__552\ : InMux
    port map (
            O => \N__4986\,
            I => \N__4983\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__4983\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_31\
        );

    \I__550\ : InMux
    port map (
            O => \N__4980\,
            I => \N__4977\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4977\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_32\
        );

    \I__548\ : InMux
    port map (
            O => \N__4974\,
            I => \N__4971\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4971\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_42\
        );

    \I__546\ : InMux
    port map (
            O => \N__4968\,
            I => \N__4965\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__4965\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_17\
        );

    \I__544\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4959\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4959\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_18\
        );

    \I__542\ : InMux
    port map (
            O => \N__4956\,
            I => \N__4953\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__4953\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_50\
        );

    \I__540\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4947\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__4947\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_51\
        );

    \I__538\ : CascadeMux
    port map (
            O => \N__4944\,
            I => \N__4940\
        );

    \I__537\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4935\
        );

    \I__536\ : InMux
    port map (
            O => \N__4940\,
            I => \N__4935\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4935\,
            I => \switch_clk_2MHz_inst.aux_CLKZ0\
        );

    \I__534\ : InMux
    port map (
            O => \N__4932\,
            I => \N__4929\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__4929\,
            I => \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_0\
        );

    \I__532\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4923\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__4923\,
            I => \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_1\
        );

    \I__530\ : InMux
    port map (
            O => \N__4920\,
            I => \N__4917\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__4917\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_8\
        );

    \I__528\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4911\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4911\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_21\
        );

    \I__526\ : InMux
    port map (
            O => \N__4908\,
            I => \N__4905\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__4905\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_66\
        );

    \I__524\ : InMux
    port map (
            O => \N__4902\,
            I => \N__4899\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4899\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_67\
        );

    \I__522\ : InMux
    port map (
            O => \N__4896\,
            I => \N__4893\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4893\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_30\
        );

    \I__520\ : InMux
    port map (
            O => \N__4890\,
            I => \N__4887\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__4887\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_28\
        );

    \I__518\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4881\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4881\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_29\
        );

    \I__516\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4875\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4875\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_38\
        );

    \I__514\ : InMux
    port map (
            O => \N__4872\,
            I => \N__4869\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4869\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_20\
        );

    \I__512\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4863\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__4863\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_19\
        );

    \I__510\ : InMux
    port map (
            O => \N__4860\,
            I => \N__4857\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4857\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_0\
        );

    \I__508\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4851\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__4851\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_1\
        );

    \I__506\ : InMux
    port map (
            O => \N__4848\,
            I => \N__4845\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4845\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_3\
        );

    \I__504\ : InMux
    port map (
            O => \N__4842\,
            I => \N__4839\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4839\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_4\
        );

    \I__502\ : InMux
    port map (
            O => \N__4836\,
            I => \N__4833\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__4833\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_5\
        );

    \I__500\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4827\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4827\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_68\
        );

    \I__498\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4821\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4821\,
            I => \N__4818\
        );

    \I__496\ : Odrv4
    port map (
            O => \N__4818\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_80\
        );

    \I__495\ : InMux
    port map (
            O => \N__4815\,
            I => \N__4812\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4812\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_64\
        );

    \I__493\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4806\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__4806\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_65\
        );

    \I__491\ : InMux
    port map (
            O => \N__4803\,
            I => \N__4800\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4800\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_12\
        );

    \I__489\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4794\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4794\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_9\
        );

    \I__487\ : InMux
    port map (
            O => \N__4791\,
            I => \N__4788\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__4788\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_10\
        );

    \I__485\ : InMux
    port map (
            O => \N__4785\,
            I => \N__4782\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4782\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_11\
        );

    \I__483\ : CEMux
    port map (
            O => \N__4779\,
            I => \N__4774\
        );

    \I__482\ : CEMux
    port map (
            O => \N__4778\,
            I => \N__4771\
        );

    \I__481\ : CEMux
    port map (
            O => \N__4777\,
            I => \N__4768\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__4774\,
            I => \switch_clk_2MHz_inst.current_state_fast_RNIJRTPZ0Z_1\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4771\,
            I => \switch_clk_2MHz_inst.current_state_fast_RNIJRTPZ0Z_1\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__4768\,
            I => \switch_clk_2MHz_inst.current_state_fast_RNIJRTPZ0Z_1\
        );

    \I__477\ : InMux
    port map (
            O => \N__4761\,
            I => \N__4758\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4758\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_6\
        );

    \I__475\ : InMux
    port map (
            O => \N__4755\,
            I => \N__4752\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4752\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_2\
        );

    \I__473\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4746\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4746\,
            I => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_7\
        );

    \I__471\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4740\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4740\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_0\
        );

    \I__469\ : InMux
    port map (
            O => \N__4737\,
            I => \N__4734\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4734\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_1\
        );

    \I__467\ : InMux
    port map (
            O => \N__4731\,
            I => \N__4728\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4728\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_2\
        );

    \I__465\ : InMux
    port map (
            O => \N__4725\,
            I => \N__4722\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4722\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_3\
        );

    \I__463\ : InMux
    port map (
            O => \N__4719\,
            I => \N__4716\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__4716\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_4\
        );

    \I__461\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4710\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__4710\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_13\
        );

    \I__459\ : InMux
    port map (
            O => \N__4707\,
            I => \N__4704\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4704\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_14\
        );

    \I__457\ : InMux
    port map (
            O => \N__4701\,
            I => \N__4698\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__4698\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_35\
        );

    \I__455\ : InMux
    port map (
            O => \N__4695\,
            I => \N__4692\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__4692\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_34\
        );

    \I__453\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4686\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4686\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_37\
        );

    \I__451\ : InMux
    port map (
            O => \N__4683\,
            I => \N__4680\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4680\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_43\
        );

    \I__449\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4674\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4674\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_52\
        );

    \I__447\ : InMux
    port map (
            O => \N__4671\,
            I => \N__4668\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__4668\,
            I => \N__4665\
        );

    \I__445\ : Odrv4
    port map (
            O => \N__4665\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_74\
        );

    \I__444\ : InMux
    port map (
            O => \N__4662\,
            I => \N__4659\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__4659\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_75\
        );

    \I__442\ : InMux
    port map (
            O => \N__4656\,
            I => \N__4653\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__4653\,
            I => \N__4650\
        );

    \I__440\ : Odrv4
    port map (
            O => \N__4650\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_16\
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__4647\,
            I => \switch_clk_2MHz_inst.counter_idlelde_2_cascade_\
        );

    \I__438\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4641\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__4641\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_15\
        );

    \I__436\ : InMux
    port map (
            O => \N__4638\,
            I => \N__4635\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__4635\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_73\
        );

    \I__434\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4629\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__4629\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_9\
        );

    \I__432\ : InMux
    port map (
            O => \N__4626\,
            I => \N__4623\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__4623\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_56\
        );

    \I__430\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4617\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__4617\,
            I => \N__4614\
        );

    \I__428\ : Odrv4
    port map (
            O => \N__4614\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_57\
        );

    \I__427\ : InMux
    port map (
            O => \N__4611\,
            I => \N__4608\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__4608\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_27\
        );

    \I__425\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4602\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__4602\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_44\
        );

    \I__423\ : InMux
    port map (
            O => \N__4599\,
            I => \N__4596\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__4596\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_26\
        );

    \I__421\ : InMux
    port map (
            O => \N__4593\,
            I => \N__4590\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__4590\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_5\
        );

    \I__419\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4584\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__4584\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_6\
        );

    \I__417\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4578\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__4578\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_7\
        );

    \I__415\ : InMux
    port map (
            O => \N__4575\,
            I => \N__4572\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__4572\,
            I => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_8\
        );

    \I__413\ : IoInMux
    port map (
            O => \N__4569\,
            I => \N__4566\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__4566\,
            I => \N__4563\
        );

    \I__411\ : IoSpan4Mux
    port map (
            O => \N__4563\,
            I => \N__4560\
        );

    \I__410\ : IoSpan4Mux
    port map (
            O => \N__4560\,
            I => \N__4557\
        );

    \I__409\ : Odrv4
    port map (
            O => \N__4557\,
            I => \RST_N_c_i\
        );

    \I__408\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4551\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__4551\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_14\
        );

    \I__406\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4545\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__4545\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_78\
        );

    \I__404\ : InMux
    port map (
            O => \N__4542\,
            I => \N__4539\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__4539\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_10\
        );

    \I__402\ : InMux
    port map (
            O => \N__4536\,
            I => \N__4533\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__4533\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_55\
        );

    \I__400\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4527\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__4527\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_76\
        );

    \I__398\ : InMux
    port map (
            O => \N__4524\,
            I => \N__4521\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__4521\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_77\
        );

    \I__396\ : InMux
    port map (
            O => \N__4518\,
            I => \N__4515\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__4515\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_36\
        );

    \I__394\ : InMux
    port map (
            O => \N__4512\,
            I => \N__4509\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__4509\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_53\
        );

    \I__392\ : InMux
    port map (
            O => \N__4506\,
            I => \N__4503\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__4503\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_54\
        );

    \I__390\ : InMux
    port map (
            O => \N__4500\,
            I => \N__4497\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__4497\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_13\
        );

    \I__388\ : InMux
    port map (
            O => \N__4494\,
            I => \N__4491\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__4491\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_12\
        );

    \I__386\ : InMux
    port map (
            O => \N__4488\,
            I => \N__4485\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__4485\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_79\
        );

    \I__384\ : InMux
    port map (
            O => \N__4482\,
            I => \N__4479\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__4479\,
            I => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_11\
        );

    \I__382\ : IoInMux
    port map (
            O => \N__4476\,
            I => \N__4473\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__4473\,
            I => \N__4470\
        );

    \I__380\ : Span12Mux_s2_v
    port map (
            O => \N__4470\,
            I => \N__4467\
        );

    \I__379\ : Span12Mux_h
    port map (
            O => \N__4467\,
            I => \N__4464\
        );

    \I__378\ : Odrv12
    port map (
            O => \N__4464\,
            I => \CLK_ibuf_gb_io_gb_input\
        );

    \IN_MUX_bfv_4_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_20_0_\
        );

    \IN_MUX_bfv_3_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_21_0_\
        );

    \IN_MUX_bfv_4_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_22_0_\
        );

    \IN_MUX_bfv_4_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_23_0_\
        );

    \CLK_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4476\,
            GLOBALBUFFEROUTPUT => \CLK_1_c_g\
        );

    \RST_N_ibuf_RNIBJGC_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4569\,
            GLOBALBUFFEROUTPUT => \RST_N_c_i_g\
        );

    \switch_clk_2MHz_inst.current_state_fast_fast_RNI0KTV_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7266\,
            GLOBALBUFFEROUTPUT => \switch_clk_2MHz_inst.N_259_g\
        );

    \switch_clk_1MHz_inst.current_state_RNITOE91_1_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6273\,
            GLOBALBUFFEROUTPUT => \switch_clk_1MHz_inst.N_377_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_13_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7980\,
            in1 => \N__6940\,
            in2 => \_gnd_net_\,
            in3 => \N__4494\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9834\,
            ce => \N__6565\,
            sr => \N__9471\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_80_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__6941\,
            in1 => \N__4488\,
            in2 => \_gnd_net_\,
            in3 => \N__7983\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9834\,
            ce => \N__6565\,
            sr => \N__9471\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_14_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5904\,
            in1 => \N__4500\,
            in2 => \_gnd_net_\,
            in3 => \N__7982\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9834\,
            ce => \N__6565\,
            sr => \N__9471\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_12_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5903\,
            in1 => \N__4482\,
            in2 => \_gnd_net_\,
            in3 => \N__7981\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9834\,
            ce => \N__6565\,
            sr => \N__9471\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_55_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__4506\,
            in1 => \N__6935\,
            in2 => \_gnd_net_\,
            in3 => \N__7995\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9832\,
            ce => \N__6567\,
            sr => \N__9472\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_79_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7992\,
            in1 => \N__6757\,
            in2 => \_gnd_net_\,
            in3 => \N__4548\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9832\,
            ce => \N__6567\,
            sr => \N__9472\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_11_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5882\,
            in1 => \N__4542\,
            in2 => \_gnd_net_\,
            in3 => \N__7994\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9832\,
            ce => \N__6567\,
            sr => \N__9472\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_78_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7991\,
            in1 => \N__6756\,
            in2 => \_gnd_net_\,
            in3 => \N__4524\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9832\,
            ce => \N__6567\,
            sr => \N__9472\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_10_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5881\,
            in1 => \N__4632\,
            in2 => \_gnd_net_\,
            in3 => \N__7993\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9832\,
            ce => \N__6567\,
            sr => \N__9472\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_56_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7990\,
            in2 => \N__6945\,
            in3 => \N__4536\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9832\,
            ce => \N__6567\,
            sr => \N__9472\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_36_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__6738\,
            in1 => \N__4701\,
            in2 => \_gnd_net_\,
            in3 => \N__7862\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9829\,
            ce => \N__6569\,
            sr => \N__9474\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_76_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7861\,
            in1 => \N__6744\,
            in2 => \_gnd_net_\,
            in3 => \N__4662\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9829\,
            ce => \N__6569\,
            sr => \N__9474\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_53_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101010101111"
        )
    port map (
            in0 => \N__4677\,
            in1 => \_gnd_net_\,
            in2 => \N__6758\,
            in3 => \N__7863\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9829\,
            ce => \N__6569\,
            sr => \N__9474\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_77_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__6927\,
            in1 => \N__4530\,
            in2 => \_gnd_net_\,
            in3 => \N__7865\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9829\,
            ce => \N__6569\,
            sr => \N__9474\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_37_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7860\,
            in1 => \N__6739\,
            in2 => \_gnd_net_\,
            in3 => \N__4518\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9829\,
            ce => \N__6569\,
            sr => \N__9474\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_54_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__6743\,
            in1 => \N__4512\,
            in2 => \_gnd_net_\,
            in3 => \N__7864\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9829\,
            ce => \N__6569\,
            sr => \N__9474\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_5_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__5889\,
            in1 => \N__4719\,
            in2 => \_gnd_net_\,
            in3 => \N__7911\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9825\,
            ce => \N__4778\,
            sr => \N__9477\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_6_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7909\,
            in1 => \N__5890\,
            in2 => \_gnd_net_\,
            in3 => \N__4593\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9825\,
            ce => \N__4778\,
            sr => \N__9477\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_7_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5891\,
            in1 => \N__4587\,
            in2 => \_gnd_net_\,
            in3 => \N__7912\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9825\,
            ce => \N__4778\,
            sr => \N__9477\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_9_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__5893\,
            in1 => \N__4575\,
            in2 => \_gnd_net_\,
            in3 => \N__7913\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9825\,
            ce => \N__4778\,
            sr => \N__9477\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_8_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7910\,
            in1 => \N__5892\,
            in2 => \_gnd_net_\,
            in3 => \N__4581\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9825\,
            ce => \N__4778\,
            sr => \N__9477\
        );

    \RST_N_ibuf_RNIBJGC_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8781\,
            lcout => \RST_N_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_58_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__6943\,
            in1 => \N__4620\,
            in2 => \_gnd_net_\,
            in3 => \N__7988\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9833\,
            ce => \N__6566\,
            sr => \N__9473\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_74_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7986\,
            in1 => \N__6755\,
            in2 => \_gnd_net_\,
            in3 => \N__4638\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9833\,
            ce => \N__6566\,
            sr => \N__9473\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_15_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5902\,
            in1 => \N__4554\,
            in2 => \_gnd_net_\,
            in3 => \N__7987\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9833\,
            ce => \N__6566\,
            sr => \N__9473\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_16_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7984\,
            in1 => \N__6942\,
            in2 => \_gnd_net_\,
            in3 => \N__4644\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9833\,
            ce => \N__6566\,
            sr => \N__9473\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_69_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__6754\,
            in1 => \N__4830\,
            in2 => \_gnd_net_\,
            in3 => \N__7989\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9833\,
            ce => \N__6566\,
            sr => \N__9473\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_73_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__7985\,
            in1 => \N__5049\,
            in2 => \_gnd_net_\,
            in3 => \N__6944\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9833\,
            ce => \N__6566\,
            sr => \N__9473\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_44_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110101111101011"
        )
    port map (
            in0 => \N__4683\,
            in1 => \N__6750\,
            in2 => \N__7972\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9830\,
            ce => \N__6570\,
            sr => \N__9475\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_28_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7894\,
            in2 => \N__6759\,
            in3 => \N__4611\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9830\,
            ce => \N__6570\,
            sr => \N__9475\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_9_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110110111101101"
        )
    port map (
            in0 => \N__6934\,
            in1 => \N__4920\,
            in2 => \N__7973\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9830\,
            ce => \N__6570\,
            sr => \N__9475\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_57_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7908\,
            in1 => \N__6933\,
            in2 => \_gnd_net_\,
            in3 => \N__4626\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9830\,
            ce => \N__6570\,
            sr => \N__9475\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_27_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100100001001000"
        )
    port map (
            in0 => \N__5880\,
            in1 => \N__4599\,
            in2 => \N__7971\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9830\,
            ce => \N__6570\,
            sr => \N__9475\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_45_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7907\,
            in1 => \N__6932\,
            in2 => \_gnd_net_\,
            in3 => \N__4605\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9830\,
            ce => \N__6570\,
            sr => \N__9475\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_26_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100100001001000"
        )
    port map (
            in0 => \N__5879\,
            in1 => \N__5193\,
            in2 => \N__7970\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9830\,
            ce => \N__6570\,
            sr => \N__9475\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_35_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__6924\,
            in1 => \N__4695\,
            in2 => \_gnd_net_\,
            in3 => \N__7878\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9826\,
            ce => \N__6572\,
            sr => \N__9478\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_34_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7874\,
            in1 => \N__6923\,
            in2 => \_gnd_net_\,
            in3 => \N__4992\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9826\,
            ce => \N__6572\,
            sr => \N__9478\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_38_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__6925\,
            in1 => \N__4689\,
            in2 => \_gnd_net_\,
            in3 => \N__7879\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9826\,
            ce => \N__6572\,
            sr => \N__9478\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_43_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7875\,
            in1 => \N__6926\,
            in2 => \_gnd_net_\,
            in3 => \N__4974\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9826\,
            ce => \N__6572\,
            sr => \N__9478\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_52_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__6736\,
            in1 => \N__4950\,
            in2 => \_gnd_net_\,
            in3 => \N__7880\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9826\,
            ce => \N__6572\,
            sr => \N__9478\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_75_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7876\,
            in1 => \N__6737\,
            in2 => \_gnd_net_\,
            in3 => \N__4671\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9826\,
            ce => \N__6572\,
            sr => \N__9478\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_17_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__4656\,
            in1 => \N__5875\,
            in2 => \_gnd_net_\,
            in3 => \N__7877\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9826\,
            ce => \N__6572\,
            sr => \N__9478\
        );

    \switch_clk_2MHz_inst.counter_idle_RNIQLMJ_5_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5474\,
            in1 => \N__5456\,
            in2 => \N__5241\,
            in3 => \N__5260\,
            lcout => OPEN,
            ltout => \switch_clk_2MHz_inst.counter_idlelde_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.current_state_fast_RNIDHKD1_1_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__7914\,
            in1 => \N__6237\,
            in2 => \N__4647\,
            in3 => \N__7416\,
            lcout => \switch_clk_2MHz_inst.current_state_fast_RNIDHKD1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.current_state_fast_RNIJRTP_1_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__7417\,
            in1 => \N__6233\,
            in2 => \_gnd_net_\,
            in3 => \N__7915\,
            lcout => \switch_clk_2MHz_inst.current_state_fast_RNIJRTPZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_0_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__7916\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6238\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9821\,
            ce => \N__4777\,
            sr => \N__9481\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_1_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__4743\,
            in1 => \N__6234\,
            in2 => \_gnd_net_\,
            in3 => \N__7919\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9821\,
            ce => \N__4777\,
            sr => \N__9481\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_2_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__7917\,
            in1 => \N__4737\,
            in2 => \_gnd_net_\,
            in3 => \N__6239\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9821\,
            ce => \N__4777\,
            sr => \N__9481\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_3_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__4731\,
            in1 => \N__6235\,
            in2 => \_gnd_net_\,
            in3 => \N__7920\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9821\,
            ce => \N__4777\,
            sr => \N__9481\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_4_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__7918\,
            in1 => \N__4725\,
            in2 => \_gnd_net_\,
            in3 => \N__6240\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9821\,
            ce => \N__4777\,
            sr => \N__9481\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_13_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5886\,
            in1 => \N__4803\,
            in2 => \_gnd_net_\,
            in3 => \N__7978\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9817\,
            ce => \N__4779\,
            sr => \N__9485\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_14_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7975\,
            in1 => \N__5887\,
            in2 => \_gnd_net_\,
            in3 => \N__4713\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9817\,
            ce => \N__4779\,
            sr => \N__9485\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_15_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5888\,
            in1 => \N__4707\,
            in2 => \_gnd_net_\,
            in3 => \N__7979\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9817\,
            ce => \N__4779\,
            sr => \N__9485\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_12_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7974\,
            in1 => \N__5885\,
            in2 => \_gnd_net_\,
            in3 => \N__4785\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9817\,
            ce => \N__4779\,
            sr => \N__9485\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_10_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5883\,
            in1 => \N__4797\,
            in2 => \_gnd_net_\,
            in3 => \N__7976\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9817\,
            ce => \N__4779\,
            sr => \N__9485\
        );

    \switch_clk_2MHz_inst.bit_sequence_din_11_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5884\,
            in1 => \N__4791\,
            in2 => \_gnd_net_\,
            in3 => \N__7977\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_dinZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9817\,
            ce => \N__4779\,
            sr => \N__9485\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_3_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10894\,
            in2 => \N__10381\,
            in3 => \N__4755\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9812\,
            ce => \N__5067\,
            sr => \N__9489\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_6_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10895\,
            in2 => \N__10382\,
            in3 => \N__4836\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9812\,
            ce => \N__5067\,
            sr => \N__9489\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_0_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__10898\,
            in1 => \N__10295\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9812\,
            ce => \N__5067\,
            sr => \N__9489\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_7_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10896\,
            in2 => \N__10383\,
            in3 => \N__4761\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9812\,
            ce => \N__5067\,
            sr => \N__9489\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_2_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110101111101011"
        )
    port map (
            in0 => \N__4854\,
            in1 => \N__10309\,
            in2 => \N__10964\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9812\,
            ce => \N__5067\,
            sr => \N__9489\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_8_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10897\,
            in2 => \N__10384\,
            in3 => \N__4749\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9812\,
            ce => \N__5067\,
            sr => \N__9489\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_1_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100000101000"
        )
    port map (
            in0 => \N__4860\,
            in1 => \N__10308\,
            in2 => \N__10963\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9812\,
            ce => \N__5067\,
            sr => \N__9489\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_4_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__4848\,
            in1 => \_gnd_net_\,
            in2 => \N__10408\,
            in3 => \N__10893\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9808\,
            ce => \N__5065\,
            sr => \N__9494\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_5_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__10892\,
            in1 => \N__10343\,
            in2 => \_gnd_net_\,
            in3 => \N__4842\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9808\,
            ce => \N__5065\,
            sr => \N__9494\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_64_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7881\,
            in1 => \N__6939\,
            in2 => \_gnd_net_\,
            in3 => \N__5127\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9831\,
            ce => \N__6568\,
            sr => \N__9476\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_22_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5878\,
            in1 => \N__4914\,
            in2 => \_gnd_net_\,
            in3 => \N__7884\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9831\,
            ce => \N__6568\,
            sr => \N__9476\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_68_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7883\,
            in1 => \N__6752\,
            in2 => \_gnd_net_\,
            in3 => \N__4902\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9831\,
            ce => \N__6568\,
            sr => \N__9476\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_81_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__6753\,
            in1 => \N__4824\,
            in2 => \_gnd_net_\,
            in3 => \N__7885\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9831\,
            ce => \N__6568\,
            sr => \N__9476\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_65_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7882\,
            in1 => \N__6751\,
            in2 => \_gnd_net_\,
            in3 => \N__4815\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9831\,
            ce => \N__6568\,
            sr => \N__9476\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_66_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7887\,
            in1 => \N__6930\,
            in2 => \_gnd_net_\,
            in3 => \N__4809\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9827\,
            ce => \N__6573\,
            sr => \N__9479\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_31_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__6929\,
            in1 => \N__4896\,
            in2 => \_gnd_net_\,
            in3 => \N__7893\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9827\,
            ce => \N__6573\,
            sr => \N__9479\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_8_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7889\,
            in1 => \N__6931\,
            in2 => \_gnd_net_\,
            in3 => \N__5205\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9827\,
            ce => \N__6573\,
            sr => \N__9479\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_21_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5876\,
            in1 => \N__4872\,
            in2 => \_gnd_net_\,
            in3 => \N__7890\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9827\,
            ce => \N__6573\,
            sr => \N__9479\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_67_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7888\,
            in1 => \N__6746\,
            in2 => \_gnd_net_\,
            in3 => \N__4908\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9827\,
            ce => \N__6573\,
            sr => \N__9479\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_30_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__6928\,
            in1 => \N__4884\,
            in2 => \_gnd_net_\,
            in3 => \N__7892\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9827\,
            ce => \N__6573\,
            sr => \N__9479\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_50_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7886\,
            in1 => \N__6745\,
            in2 => \_gnd_net_\,
            in3 => \N__5220\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9827\,
            ce => \N__6573\,
            sr => \N__9479\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_29_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5877\,
            in1 => \N__4890\,
            in2 => \_gnd_net_\,
            in3 => \N__7891\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9827\,
            ce => \N__6573\,
            sr => \N__9479\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_39_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__6921\,
            in1 => \N__4878\,
            in2 => \_gnd_net_\,
            in3 => \N__7873\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9822\,
            ce => \N__6575\,
            sr => \N__9482\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_20_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7866\,
            in1 => \N__5874\,
            in2 => \_gnd_net_\,
            in3 => \N__4866\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9822\,
            ce => \N__6575\,
            sr => \N__9482\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_19_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5873\,
            in1 => \N__4962\,
            in2 => \_gnd_net_\,
            in3 => \N__7871\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9822\,
            ce => \N__6575\,
            sr => \N__9482\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_33_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7867\,
            in1 => \N__6684\,
            in2 => \_gnd_net_\,
            in3 => \N__4980\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9822\,
            ce => \N__6575\,
            sr => \N__9482\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_32_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__6920\,
            in1 => \N__4986\,
            in2 => \_gnd_net_\,
            in3 => \N__7872\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9822\,
            ce => \N__6575\,
            sr => \N__9482\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_42_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7868\,
            in1 => \N__6685\,
            in2 => \_gnd_net_\,
            in3 => \N__6963\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9822\,
            ce => \N__6575\,
            sr => \N__9482\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_18_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5872\,
            in1 => \N__4968\,
            in2 => \_gnd_net_\,
            in3 => \N__7870\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9822\,
            ce => \N__6575\,
            sr => \N__9482\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_51_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7869\,
            in1 => \N__6922\,
            in2 => \_gnd_net_\,
            in3 => \N__4956\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9822\,
            ce => \N__6575\,
            sr => \N__9482\
        );

    \switch_clk_2MHz_inst.delay_inst.delay_reg_1_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4932\,
            lcout => \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9818\,
            ce => 'H',
            sr => \N__9486\
        );

    \switch_clk_2MHz_inst.aux_CLK_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011010010000"
        )
    port map (
            in0 => \N__7808\,
            in1 => \N__6236\,
            in2 => \N__4944\,
            in3 => \N__7299\,
            lcout => \switch_clk_2MHz_inst.aux_CLKZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9818\,
            ce => 'H',
            sr => \N__9486\
        );

    \switch_clk_2MHz_inst.delay_inst.delay_reg_0_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4943\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9818\,
            ce => 'H',
            sr => \N__9486\
        );

    \switch_clk_2MHz_inst.delay_inst.delay_reg_2_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4926\,
            lcout => \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9818\,
            ce => 'H',
            sr => \N__9486\
        );

    \switch_clk_2MHz_inst.counter_idle_0_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5425\,
            in1 => \N__5286\,
            in2 => \_gnd_net_\,
            in3 => \N__5034\,
            lcout => \switch_clk_2MHz_inst.counter_idleZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_21_0_\,
            carryout => \switch_clk_2MHz_inst.counter_idle_cry_0\,
            clk => \N__9813\,
            ce => \N__5016\,
            sr => \N__9490\
        );

    \switch_clk_2MHz_inst.counter_idle_1_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5422\,
            in1 => \N__5274\,
            in2 => \_gnd_net_\,
            in3 => \N__5031\,
            lcout => \switch_clk_2MHz_inst.counter_idleZ0Z_1\,
            ltout => OPEN,
            carryin => \switch_clk_2MHz_inst.counter_idle_cry_0\,
            carryout => \switch_clk_2MHz_inst.counter_idle_cry_1\,
            clk => \N__9813\,
            ce => \N__5016\,
            sr => \N__9490\
        );

    \switch_clk_2MHz_inst.counter_idle_2_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5426\,
            in1 => \N__5261\,
            in2 => \_gnd_net_\,
            in3 => \N__5028\,
            lcout => \switch_clk_2MHz_inst.counter_idleZ0Z_2\,
            ltout => OPEN,
            carryin => \switch_clk_2MHz_inst.counter_idle_cry_1\,
            carryout => \switch_clk_2MHz_inst.counter_idle_cry_2\,
            clk => \N__9813\,
            ce => \N__5016\,
            sr => \N__9490\
        );

    \switch_clk_2MHz_inst.counter_idle_3_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5423\,
            in1 => \N__5457\,
            in2 => \_gnd_net_\,
            in3 => \N__5025\,
            lcout => \switch_clk_2MHz_inst.counter_idleZ0Z_3\,
            ltout => OPEN,
            carryin => \switch_clk_2MHz_inst.counter_idle_cry_2\,
            carryout => \switch_clk_2MHz_inst.counter_idle_cry_3\,
            clk => \N__9813\,
            ce => \N__5016\,
            sr => \N__9490\
        );

    \switch_clk_2MHz_inst.counter_idle_4_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5427\,
            in1 => \N__5475\,
            in2 => \_gnd_net_\,
            in3 => \N__5022\,
            lcout => \switch_clk_2MHz_inst.counter_idleZ0Z_4\,
            ltout => OPEN,
            carryin => \switch_clk_2MHz_inst.counter_idle_cry_3\,
            carryout => \switch_clk_2MHz_inst.counter_idle_cry_4\,
            clk => \N__9813\,
            ce => \N__5016\,
            sr => \N__9490\
        );

    \switch_clk_2MHz_inst.counter_idle_5_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5424\,
            in1 => \N__5240\,
            in2 => \_gnd_net_\,
            in3 => \N__5019\,
            lcout => \switch_clk_2MHz_inst.counter_idleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9813\,
            ce => \N__5016\,
            sr => \N__9490\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_10_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__4998\,
            in1 => \_gnd_net_\,
            in2 => \N__10347\,
            in3 => \N__10764\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9809\,
            ce => \N__5066\,
            sr => \N__9495\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_9_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__10763\,
            in1 => \N__10229\,
            in2 => \_gnd_net_\,
            in3 => \N__5004\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9809\,
            ce => \N__5066\,
            sr => \N__9495\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_12_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__5094\,
            in1 => \_gnd_net_\,
            in2 => \N__10349\,
            in3 => \N__10766\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9809\,
            ce => \N__5066\,
            sr => \N__9495\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_15_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__10762\,
            in1 => \N__10228\,
            in2 => \_gnd_net_\,
            in3 => \N__5088\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9809\,
            ce => \N__5066\,
            sr => \N__9495\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_11_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101010101111"
        )
    port map (
            in0 => \N__5100\,
            in1 => \_gnd_net_\,
            in2 => \N__10348\,
            in3 => \N__10765\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9809\,
            ce => \N__5066\,
            sr => \N__9495\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_14_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__10761\,
            in1 => \N__10227\,
            in2 => \_gnd_net_\,
            in3 => \N__5076\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9809\,
            ce => \N__5066\,
            sr => \N__9495\
        );

    \switch_clk_1MHz_inst.bit_sequence_din_13_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101010101111"
        )
    port map (
            in0 => \N__5082\,
            in1 => \_gnd_net_\,
            in2 => \N__10350\,
            in3 => \N__10767\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_dinZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9809\,
            ce => \N__5066\,
            sr => \N__9495\
        );

    \switch_clk_1MHz_inst.counter_stat_RNIIHP11_6_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__5971\,
            in1 => \N__5369\,
            in2 => \N__5531\,
            in3 => \N__6002\,
            lcout => OPEN,
            ltout => \switch_clk_1MHz_inst.counter_statlde_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_RNIFA8B2_1_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100000000"
        )
    port map (
            in0 => \N__10759\,
            in1 => \N__9979\,
            in2 => \N__5070\,
            in3 => \N__9089\,
            lcout => \switch_clk_1MHz_inst.current_state_RNIFA8B2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_RNITOE91_1_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__9090\,
            in1 => \N__10760\,
            in2 => \_gnd_net_\,
            in3 => \N__9998\,
            lcout => \switch_clk_1MHz_inst.current_state_RNITOE91Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_72_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7825\,
            in1 => \N__6883\,
            in2 => \_gnd_net_\,
            in3 => \N__5145\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9828\,
            ce => \N__6571\,
            sr => \N__9480\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_82_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__6729\,
            in1 => \N__5040\,
            in2 => \_gnd_net_\,
            in3 => \N__7829\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9828\,
            ce => \N__6571\,
            sr => \N__9480\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_70_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7824\,
            in1 => \N__6882\,
            in2 => \_gnd_net_\,
            in3 => \N__5160\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9828\,
            ce => \N__6571\,
            sr => \N__9480\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_71_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__6728\,
            in1 => \N__5151\,
            in2 => \_gnd_net_\,
            in3 => \N__7828\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9828\,
            ce => \N__6571\,
            sr => \N__9480\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_23_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7822\,
            in1 => \N__5832\,
            in2 => \_gnd_net_\,
            in3 => \N__5139\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9828\,
            ce => \N__6571\,
            sr => \N__9480\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_62_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__6881\,
            in1 => \N__5676\,
            in2 => \_gnd_net_\,
            in3 => \N__7827\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9828\,
            ce => \N__6571\,
            sr => \N__9480\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_63_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7823\,
            in1 => \N__6727\,
            in2 => \_gnd_net_\,
            in3 => \N__5133\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9828\,
            ce => \N__6571\,
            sr => \N__9480\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_59_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__6726\,
            in1 => \N__5121\,
            in2 => \_gnd_net_\,
            in3 => \N__7826\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9828\,
            ce => \N__6571\,
            sr => \N__9480\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_24_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5792\,
            in1 => \N__5112\,
            in2 => \_gnd_net_\,
            in3 => \N__7818\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9823\,
            ce => \N__6576\,
            sr => \N__9483\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_5_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7816\,
            in1 => \N__5796\,
            in2 => \_gnd_net_\,
            in3 => \N__5106\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9823\,
            ce => \N__6576\,
            sr => \N__9483\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_4_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5795\,
            in1 => \N__5184\,
            in2 => \_gnd_net_\,
            in3 => \N__7821\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9823\,
            ce => \N__6576\,
            sr => \N__9483\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_49_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7815\,
            in1 => \N__6675\,
            in2 => \_gnd_net_\,
            in3 => \N__5925\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9823\,
            ce => \N__6576\,
            sr => \N__9483\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_46_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__6674\,
            in1 => \N__5214\,
            in2 => \_gnd_net_\,
            in3 => \N__7820\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9823\,
            ce => \N__6576\,
            sr => \N__9483\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_7_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__7817\,
            in1 => \_gnd_net_\,
            in2 => \N__5343\,
            in3 => \N__5797\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9823\,
            ce => \N__6576\,
            sr => \N__9483\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_25_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__5793\,
            in1 => \N__5199\,
            in2 => \_gnd_net_\,
            in3 => \N__7819\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9823\,
            ce => \N__6576\,
            sr => \N__9483\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_3_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7814\,
            in1 => \N__5794\,
            in2 => \_gnd_net_\,
            in3 => \N__5166\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9823\,
            ce => \N__6576\,
            sr => \N__9483\
        );

    \switch_clk_2MHz_inst.current_state_RNO_0_0_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7462\,
            in1 => \N__5334\,
            in2 => \N__5316\,
            in3 => \N__6257\,
            lcout => \switch_clk_2MHz_inst.G_31_0_a4_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_0_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7463\,
            in2 => \_gnd_net_\,
            in3 => \N__7689\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9819\,
            ce => \N__6577\,
            sr => \N__9487\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_1_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7688\,
            in1 => \N__5777\,
            in2 => \_gnd_net_\,
            in3 => \N__5178\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9819\,
            ce => \N__6577\,
            sr => \N__9487\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_2_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__6818\,
            in1 => \N__5172\,
            in2 => \_gnd_net_\,
            in3 => \N__7690\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9819\,
            ce => \N__6577\,
            sr => \N__9487\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_6_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__6819\,
            in1 => \N__5349\,
            in2 => \_gnd_net_\,
            in3 => \N__7691\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9819\,
            ce => \N__6577\,
            sr => \N__9487\
        );

    \switch_clk_2MHz_inst.counter_stat_0_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5728\,
            in1 => \N__5333\,
            in2 => \_gnd_net_\,
            in3 => \N__5322\,
            lcout => \switch_clk_2MHz_inst.counter_statZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_20_0_\,
            carryout => \switch_clk_2MHz_inst.counter_stat_cry_0\,
            clk => \N__9814\,
            ce => \N__6180\,
            sr => \N__9491\
        );

    \switch_clk_2MHz_inst.counter_stat_1_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5724\,
            in1 => \N__6171\,
            in2 => \_gnd_net_\,
            in3 => \N__5319\,
            lcout => \switch_clk_2MHz_inst.counter_statZ0Z_1\,
            ltout => OPEN,
            carryin => \switch_clk_2MHz_inst.counter_stat_cry_0\,
            carryout => \switch_clk_2MHz_inst.counter_stat_cry_1\,
            clk => \N__9814\,
            ce => \N__6180\,
            sr => \N__9491\
        );

    \switch_clk_2MHz_inst.counter_stat_2_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5729\,
            in1 => \N__5312\,
            in2 => \_gnd_net_\,
            in3 => \N__5301\,
            lcout => \switch_clk_2MHz_inst.counter_statZ0Z_2\,
            ltout => OPEN,
            carryin => \switch_clk_2MHz_inst.counter_stat_cry_1\,
            carryout => \switch_clk_2MHz_inst.counter_stat_cry_2\,
            clk => \N__9814\,
            ce => \N__6180\,
            sr => \N__9491\
        );

    \switch_clk_2MHz_inst.counter_stat_3_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5725\,
            in1 => \N__6258\,
            in2 => \_gnd_net_\,
            in3 => \N__5298\,
            lcout => \switch_clk_2MHz_inst.counter_statZ0Z_3\,
            ltout => OPEN,
            carryin => \switch_clk_2MHz_inst.counter_stat_cry_2\,
            carryout => \switch_clk_2MHz_inst.counter_stat_cry_3\,
            clk => \N__9814\,
            ce => \N__6180\,
            sr => \N__9491\
        );

    \switch_clk_2MHz_inst.counter_stat_4_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5730\,
            in1 => \N__6118\,
            in2 => \_gnd_net_\,
            in3 => \N__5295\,
            lcout => \switch_clk_2MHz_inst.counter_statZ0Z_4\,
            ltout => OPEN,
            carryin => \switch_clk_2MHz_inst.counter_stat_cry_3\,
            carryout => \switch_clk_2MHz_inst.counter_stat_cry_4\,
            clk => \N__9814\,
            ce => \N__6180\,
            sr => \N__9491\
        );

    \switch_clk_2MHz_inst.counter_stat_5_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5726\,
            in1 => \N__6139\,
            in2 => \_gnd_net_\,
            in3 => \N__5292\,
            lcout => \switch_clk_2MHz_inst.counter_statZ0Z_5\,
            ltout => OPEN,
            carryin => \switch_clk_2MHz_inst.counter_stat_cry_4\,
            carryout => \switch_clk_2MHz_inst.counter_stat_cry_5\,
            clk => \N__9814\,
            ce => \N__6180\,
            sr => \N__9491\
        );

    \switch_clk_2MHz_inst.counter_stat_6_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__6159\,
            in1 => \N__5727\,
            in2 => \_gnd_net_\,
            in3 => \N__5289\,
            lcout => \switch_clk_2MHz_inst.counter_statZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9814\,
            ce => \N__6180\,
            sr => \N__9491\
        );

    \switch_clk_2MHz_inst.current_state_RNO_6_0_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5285\,
            in1 => \N__5273\,
            in2 => \N__5262\,
            in3 => \N__5239\,
            lcout => \switch_clk_2MHz_inst.G_31_0_a4_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.current_state_RNO_7_0_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5473\,
            in1 => \N__5455\,
            in2 => \N__5919\,
            in3 => \N__7606\,
            lcout => OPEN,
            ltout => \switch_clk_2MHz_inst.G_31_0_a4_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.current_state_RNO_3_0_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7488\,
            in1 => \N__5439\,
            in2 => \N__5433\,
            in3 => \N__7419\,
            lcout => \switch_clk_2MHz_inst.N_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_RNO_6_0_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__5368\,
            in1 => \N__5384\,
            in2 => \N__5532\,
            in3 => \N__5402\,
            lcout => OPEN,
            ltout => \switch_clk_1MHz_inst.current_state_ns_0_a3_1_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_RNO_1_0_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5430\,
            in3 => \N__5952\,
            lcout => \switch_clk_1MHz_inst.current_state_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.current_state_fast_1_rep1_RNIEUV6_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7487\,
            in2 => \_gnd_net_\,
            in3 => \N__7607\,
            lcout => \switch_clk_2MHz_inst.N_117_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.counter_stat_0_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6344\,
            in1 => \N__5403\,
            in2 => \_gnd_net_\,
            in3 => \N__5391\,
            lcout => \switch_clk_1MHz_inst.counter_statZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_22_0_\,
            carryout => \switch_clk_1MHz_inst.counter_stat_cry_0\,
            clk => \N__9804\,
            ce => \N__5508\,
            sr => \N__9498\
        );

    \switch_clk_1MHz_inst.counter_stat_1_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6355\,
            in1 => \N__5985\,
            in2 => \_gnd_net_\,
            in3 => \N__5388\,
            lcout => \switch_clk_1MHz_inst.counter_statZ0Z_1\,
            ltout => OPEN,
            carryin => \switch_clk_1MHz_inst.counter_stat_cry_0\,
            carryout => \switch_clk_1MHz_inst.counter_stat_cry_1\,
            clk => \N__9804\,
            ce => \N__5508\,
            sr => \N__9498\
        );

    \switch_clk_1MHz_inst.counter_stat_2_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6345\,
            in1 => \N__5385\,
            in2 => \_gnd_net_\,
            in3 => \N__5373\,
            lcout => \switch_clk_1MHz_inst.counter_statZ0Z_2\,
            ltout => OPEN,
            carryin => \switch_clk_1MHz_inst.counter_stat_cry_1\,
            carryout => \switch_clk_1MHz_inst.counter_stat_cry_2\,
            clk => \N__9804\,
            ce => \N__5508\,
            sr => \N__9498\
        );

    \switch_clk_1MHz_inst.counter_stat_3_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6356\,
            in1 => \N__5370\,
            in2 => \_gnd_net_\,
            in3 => \N__5352\,
            lcout => \switch_clk_1MHz_inst.counter_statZ0Z_3\,
            ltout => OPEN,
            carryin => \switch_clk_1MHz_inst.counter_stat_cry_2\,
            carryout => \switch_clk_1MHz_inst.counter_stat_cry_3\,
            clk => \N__9804\,
            ce => \N__5508\,
            sr => \N__9498\
        );

    \switch_clk_1MHz_inst.counter_stat_4_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6346\,
            in1 => \N__6003\,
            in2 => \_gnd_net_\,
            in3 => \N__5541\,
            lcout => \switch_clk_1MHz_inst.counter_statZ0Z_4\,
            ltout => OPEN,
            carryin => \switch_clk_1MHz_inst.counter_stat_cry_3\,
            carryout => \switch_clk_1MHz_inst.counter_stat_cry_4\,
            clk => \N__9804\,
            ce => \N__5508\,
            sr => \N__9498\
        );

    \switch_clk_1MHz_inst.counter_stat_5_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6357\,
            in1 => \N__5972\,
            in2 => \_gnd_net_\,
            in3 => \N__5538\,
            lcout => \switch_clk_1MHz_inst.counter_statZ0Z_5\,
            ltout => OPEN,
            carryin => \switch_clk_1MHz_inst.counter_stat_cry_4\,
            carryout => \switch_clk_1MHz_inst.counter_stat_cry_5\,
            clk => \N__9804\,
            ce => \N__5508\,
            sr => \N__9498\
        );

    \switch_clk_1MHz_inst.counter_stat_6_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6347\,
            in1 => \N__5530\,
            in2 => \_gnd_net_\,
            in3 => \N__5535\,
            lcout => \switch_clk_1MHz_inst.counter_statZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9804\,
            ce => \N__5508\,
            sr => \N__9498\
        );

    \switch_clk_1MHz_inst.counter_idle_0_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6324\,
            in1 => \N__6029\,
            in2 => \_gnd_net_\,
            in3 => \N__5493\,
            lcout => \switch_clk_1MHz_inst.counter_idleZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_23_0_\,
            carryout => \switch_clk_1MHz_inst.counter_idle_cry_0\,
            clk => \N__9800\,
            ce => \N__5637\,
            sr => \N__9502\
        );

    \switch_clk_1MHz_inst.counter_idle_1_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6320\,
            in1 => \N__6068\,
            in2 => \_gnd_net_\,
            in3 => \N__5490\,
            lcout => \switch_clk_1MHz_inst.counter_idleZ0Z_1\,
            ltout => OPEN,
            carryin => \switch_clk_1MHz_inst.counter_idle_cry_0\,
            carryout => \switch_clk_1MHz_inst.counter_idle_cry_1\,
            clk => \N__9800\,
            ce => \N__5637\,
            sr => \N__9502\
        );

    \switch_clk_1MHz_inst.counter_idle_2_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6325\,
            in1 => \N__6083\,
            in2 => \_gnd_net_\,
            in3 => \N__5487\,
            lcout => \switch_clk_1MHz_inst.counter_idleZ0Z_2\,
            ltout => OPEN,
            carryin => \switch_clk_1MHz_inst.counter_idle_cry_1\,
            carryout => \switch_clk_1MHz_inst.counter_idle_cry_2\,
            clk => \N__9800\,
            ce => \N__5637\,
            sr => \N__9502\
        );

    \switch_clk_1MHz_inst.counter_idle_3_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6321\,
            in1 => \N__5631\,
            in2 => \_gnd_net_\,
            in3 => \N__5484\,
            lcout => \switch_clk_1MHz_inst.counter_idleZ0Z_3\,
            ltout => OPEN,
            carryin => \switch_clk_1MHz_inst.counter_idle_cry_2\,
            carryout => \switch_clk_1MHz_inst.counter_idle_cry_3\,
            clk => \N__9800\,
            ce => \N__5637\,
            sr => \N__9502\
        );

    \switch_clk_1MHz_inst.counter_idle_4_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6326\,
            in1 => \N__5616\,
            in2 => \_gnd_net_\,
            in3 => \N__5481\,
            lcout => \switch_clk_1MHz_inst.counter_idleZ0Z_4\,
            ltout => OPEN,
            carryin => \switch_clk_1MHz_inst.counter_idle_cry_3\,
            carryout => \switch_clk_1MHz_inst.counter_idle_cry_4\,
            clk => \N__9800\,
            ce => \N__5637\,
            sr => \N__9502\
        );

    \switch_clk_1MHz_inst.counter_idle_5_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6322\,
            in1 => \N__6050\,
            in2 => \_gnd_net_\,
            in3 => \N__5478\,
            lcout => \switch_clk_1MHz_inst.counter_idleZ0Z_5\,
            ltout => OPEN,
            carryin => \switch_clk_1MHz_inst.counter_idle_cry_4\,
            carryout => \switch_clk_1MHz_inst.counter_idle_cry_5\,
            clk => \N__9800\,
            ce => \N__5637\,
            sr => \N__9502\
        );

    \switch_clk_1MHz_inst.counter_idle_6_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6327\,
            in1 => \N__5578\,
            in2 => \_gnd_net_\,
            in3 => \N__5652\,
            lcout => \switch_clk_1MHz_inst.counter_idleZ0Z_6\,
            ltout => OPEN,
            carryin => \switch_clk_1MHz_inst.counter_idle_cry_5\,
            carryout => \switch_clk_1MHz_inst.counter_idle_cry_6\,
            clk => \N__9800\,
            ce => \N__5637\,
            sr => \N__9502\
        );

    \switch_clk_1MHz_inst.counter_idle_7_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6323\,
            in1 => \N__5599\,
            in2 => \_gnd_net_\,
            in3 => \N__5649\,
            lcout => \switch_clk_1MHz_inst.counter_idleZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9800\,
            ce => \N__5637\,
            sr => \N__9502\
        );

    \switch_clk_1MHz_inst.current_state_RNI1TCQ_2_1_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__9945\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10508\,
            lcout => \switch_clk_1MHz_inst.N_116_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.counter_idle_RNIQP3H_3_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011111"
        )
    port map (
            in0 => \N__5630\,
            in1 => \N__6049\,
            in2 => \N__5583\,
            in3 => \N__5615\,
            lcout => OPEN,
            ltout => \switch_clk_1MHz_inst.G_31_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.counter_idle_RNIOJRU1_7_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__5646\,
            in1 => \N__5600\,
            in2 => \N__5640\,
            in3 => \N__9081\,
            lcout => \switch_clk_1MHz_inst.counter_idle_RNIOJRU1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_RNO_5_0_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5629\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5614\,
            lcout => \switch_clk_1MHz_inst.current_state_RNO_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_RNO_4_0_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__9946\,
            in1 => \N__8136\,
            in2 => \N__10771\,
            in3 => \N__5601\,
            lcout => OPEN,
            ltout => \switch_clk_1MHz_inst.current_state_RNO_4Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_RNO_0_0_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__5582\,
            in1 => \N__5562\,
            in2 => \N__5556\,
            in3 => \N__6015\,
            lcout => OPEN,
            ltout => \switch_clk_1MHz_inst.N_116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_0_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011100010111011"
        )
    port map (
            in0 => \N__9947\,
            in1 => \N__6411\,
            in2 => \N__5553\,
            in3 => \N__5550\,
            lcout => \switch_clk_1MHz_inst_current_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9797\,
            ce => 'H',
            sr => \N__9506\
        );

    \switch_clk_1MHz_inst.current_state_RNI1TCQ_1_1_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10612\,
            in3 => \N__9944\,
            lcout => \switch_clk_1MHz_inst.N_90_li\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.counter_din_RNIFO9H_1_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6457\,
            in2 => \_gnd_net_\,
            in3 => \N__6432\,
            lcout => \switch_clk_1MHz_inst.N_88_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_58_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__10678\,
            in1 => \_gnd_net_\,
            in2 => \N__6516\,
            in3 => \N__10190\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9788\,
            ce => \N__9617\,
            sr => \N__9513\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_59_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10189\,
            in1 => \N__5703\,
            in2 => \_gnd_net_\,
            in3 => \N__10679\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9788\,
            ce => \N__9617\,
            sr => \N__9513\
        );

    \config_register_latched_dec_inst.DYNCNF_1_RNIP1121_0_0_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6297\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DYNCNF_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_83_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__6725\,
            in1 => \N__5682\,
            in2 => \_gnd_net_\,
            in3 => \N__7813\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9824\,
            ce => \N__6574\,
            sr => \N__9484\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_61_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7810\,
            in1 => \N__6880\,
            in2 => \_gnd_net_\,
            in3 => \N__5658\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9824\,
            ce => \N__6574\,
            sr => \N__9484\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_47_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__6878\,
            in1 => \N__5670\,
            in2 => \_gnd_net_\,
            in3 => \N__7811\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9824\,
            ce => \N__6574\,
            sr => \N__9484\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_60_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7809\,
            in1 => \N__6724\,
            in2 => \_gnd_net_\,
            in3 => \N__5664\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9824\,
            ce => \N__6574\,
            sr => \N__9484\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_48_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__6879\,
            in1 => \N__5931\,
            in2 => \_gnd_net_\,
            in3 => \N__7812\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9824\,
            ce => \N__6574\,
            sr => \N__9484\
        );

    \switch_clk_2MHz_inst.flag_input_reg_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8325\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_2MHz_inst.flag_input_regZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9820\,
            ce => 'H',
            sr => \N__9488\
        );

    \switch_clk_2MHz_inst.current_state_fast_1_rep1_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__7415\,
            in1 => \N__7465\,
            in2 => \N__7247\,
            in3 => \N__7830\,
            lcout => \switch_clk_2MHz_inst.current_state_fast_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9820\,
            ce => 'H',
            sr => \N__9488\
        );

    \switch_clk_2MHz_inst.current_state_1_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__7609\,
            in1 => \N__7235\,
            in2 => \N__6735\,
            in3 => \N__7403\,
            lcout => \switch_clk_2MHz_inst.current_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9815\,
            ce => 'H',
            sr => \N__9492\
        );

    \switch_clk_2MHz_inst.counter_din_RNI6HAE1_3_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7049\,
            in1 => \N__7077\,
            in2 => \N__7017\,
            in3 => \N__7104\,
            lcout => \switch_clk_2MHz_inst.N_114_0\,
            ltout => \switch_clk_2MHz_inst.N_114_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.current_state_1_rep1_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__7404\,
            in1 => \N__5831\,
            in2 => \N__5907\,
            in3 => \N__7611\,
            lcout => \switch_clk_2MHz_inst.current_state_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9815\,
            ce => 'H',
            sr => \N__9492\
        );

    \switch_clk_2MHz_inst.current_state_fast_1_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__7610\,
            in1 => \N__7239\,
            in2 => \N__6232\,
            in3 => \N__7406\,
            lcout => \switch_clk_2MHz_inst.current_state_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9815\,
            ce => 'H',
            sr => \N__9492\
        );

    \switch_clk_2MHz_inst.current_state_1_rep2_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__7405\,
            in1 => \N__6858\,
            in2 => \N__7246\,
            in3 => \N__7612\,
            lcout => \switch_clk_2MHz_inst.current_state_1_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9815\,
            ce => 'H',
            sr => \N__9492\
        );

    \switch_clk_2MHz_inst.current_state_fast_1_rep1_RNIEUV6_0_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7464\,
            in2 => \_gnd_net_\,
            in3 => \N__7608\,
            lcout => \switch_clk_2MHz_inst.current_state_d_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.counter_stat_RNIMHC41_6_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__6119\,
            in1 => \N__6256\,
            in2 => \N__6144\,
            in3 => \N__6157\,
            lcout => OPEN,
            ltout => \switch_clk_2MHz_inst.counter_statlde_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.current_state_fast_RNI9DAU1_1_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100000000"
        )
    port map (
            in0 => \N__6209\,
            in1 => \N__7605\,
            in2 => \N__6183\,
            in3 => \N__7387\,
            lcout => \switch_clk_2MHz_inst.current_state_fast_RNI9DAU1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.current_state_RNO_4_0_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6170\,
            in2 => \_gnd_net_\,
            in3 => \N__6158\,
            lcout => OPEN,
            ltout => \switch_clk_2MHz_inst.G_31_0_a4_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.current_state_RNO_1_0_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6143\,
            in1 => \N__6120\,
            in2 => \N__6102\,
            in3 => \N__7386\,
            lcout => OPEN,
            ltout => \switch_clk_2MHz_inst.G_31_0_a4_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.current_state_0_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__6099\,
            in1 => \N__6093\,
            in2 => \N__6087\,
            in3 => \N__6363\,
            lcout => \switch_clk_2MHz_inst.current_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9810\,
            ce => 'H',
            sr => \N__9496\
        );

    \switch_clk_1MHz_inst.current_state_RNO_3_0_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__6084\,
            in1 => \N__6069\,
            in2 => \N__6054\,
            in3 => \N__6030\,
            lcout => \switch_clk_1MHz_inst.current_state_RNO_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_RNO_7_0_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6001\,
            in1 => \N__5984\,
            in2 => \N__5973\,
            in3 => \N__10654\,
            lcout => \switch_clk_1MHz_inst.current_state_ns_0_a3_1_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.MOSI_er_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110010000100000"
        )
    port map (
            in0 => \N__7621\,
            in1 => \N__7480\,
            in2 => \N__5946\,
            in3 => \N__6954\,
            lcout => \mosi_2MHz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9805\,
            ce => \N__7385\,
            sr => \N__9499\
        );

    \switch_clk_2MHz_inst.current_state_RNO_2_0_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001100"
        )
    port map (
            in0 => \N__7110\,
            in1 => \N__7620\,
            in2 => \N__7489\,
            in3 => \N__7384\,
            lcout => \switch_clk_2MHz_inst.N_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst.STATCNF_1_RNO_0_0_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__8024\,
            in1 => \N__10105\,
            in2 => \_gnd_net_\,
            in3 => \N__9067\,
            lcout => \config_register_latched_dec_inst.STATCNF_1_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.SEL_0_er_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10108\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \aux_selection_1MHz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9801\,
            ce => \N__9101\,
            sr => \N__9503\
        );

    \switch_clk_1MHz_inst.counter_din_RNO_0_3_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6387\,
            in1 => \N__6462\,
            in2 => \_gnd_net_\,
            in3 => \N__6440\,
            lcout => \switch_clk_1MHz_inst.N_91_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_RNI1TCQ_0_1_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__10106\,
            in1 => \_gnd_net_\,
            in2 => \N__10772\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_1MHz_inst.current_state_d_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_RNI1TCQ_1_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10655\,
            in2 => \_gnd_net_\,
            in3 => \N__10107\,
            lcout => \switch_clk_1MHz_inst.N_116_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst.DYNCNF_1_RNIP1121_0_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__6285\,
            in1 => \N__8555\,
            in2 => \N__8791\,
            in3 => \N__8706\,
            lcout => \config_register_latched_dec_inst.DYNCNF_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst.DYNCNF_1_0_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__8705\,
            in1 => \N__8782\,
            in2 => \N__8556\,
            in3 => \N__6284\,
            lcout => \config_register_latched_dec_inst.DYNCNF_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9798\,
            ce => \N__7122\,
            sr => \N__9507\
        );

    \divisor_inst_2.counter_RNISR1F_2_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8234\,
            in1 => \N__8125\,
            in2 => \N__8198\,
            in3 => \N__8212\,
            lcout => \counter_RNISR1F_2\,
            ltout => \counter_RNISR1F_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_RNITOE91_0_1_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6276\,
            in3 => \N__8081\,
            lcout => \switch_clk_1MHz_inst.current_state_RNITOE91_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_RNO_0_1_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10000\,
            in1 => \N__6382\,
            in2 => \N__8061\,
            in3 => \N__6401\,
            lcout => OPEN,
            ltout => \switch_clk_1MHz_inst.current_state_cnv_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_1_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101010101010"
        )
    port map (
            in0 => \N__10634\,
            in1 => \_gnd_net_\,
            in2 => \N__6465\,
            in3 => \N__9097\,
            lcout => \switch_clk_1MHz_inst.current_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9793\,
            ce => 'H',
            sr => \N__9509\
        );

    \switch_clk_1MHz_inst.counter_din_1_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100011001100"
        )
    port map (
            in0 => \N__8083\,
            in1 => \N__6461\,
            in2 => \N__6441\,
            in3 => \N__9080\,
            lcout => \switch_clk_1MHz_inst.counter_dinZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9793\,
            ce => 'H',
            sr => \N__9509\
        );

    \switch_clk_1MHz_inst.counter_din_0_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011001000100"
        )
    port map (
            in0 => \N__9078\,
            in1 => \N__6436\,
            in2 => \_gnd_net_\,
            in3 => \N__8082\,
            lcout => \switch_clk_1MHz_inst.counter_dinZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9793\,
            ce => 'H',
            sr => \N__9509\
        );

    \switch_clk_1MHz_inst.current_state_RNO_8_0_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8056\,
            in1 => \N__6381\,
            in2 => \_gnd_net_\,
            in3 => \N__10633\,
            lcout => OPEN,
            ltout => \switch_clk_1MHz_inst.current_state_RNO_8Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.current_state_RNO_2_0_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101010101"
        )
    port map (
            in0 => \N__9077\,
            in1 => \N__6400\,
            in2 => \N__6414\,
            in3 => \N__9999\,
            lcout => \switch_clk_1MHz_inst.current_state_RNO_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.counter_din_2_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110001000100"
        )
    port map (
            in0 => \N__9079\,
            in1 => \N__6386\,
            in2 => \N__6405\,
            in3 => \N__8084\,
            lcout => \switch_clk_1MHz_inst.counter_dinZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9793\,
            ce => 'H',
            sr => \N__9509\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_25_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__10602\,
            in1 => \N__10098\,
            in2 => \_gnd_net_\,
            in3 => \N__6528\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9789\,
            ce => \N__9618\,
            sr => \N__9514\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_28_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__6501\,
            in1 => \N__10607\,
            in2 => \_gnd_net_\,
            in3 => \N__10103\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9789\,
            ce => \N__9618\,
            sr => \N__9514\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_24_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__10601\,
            in1 => \N__10097\,
            in2 => \_gnd_net_\,
            in3 => \N__6507\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9789\,
            ce => \N__9618\,
            sr => \N__9514\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_29_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__6522\,
            in1 => \N__10608\,
            in2 => \_gnd_net_\,
            in3 => \N__10104\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9789\,
            ce => \N__9618\,
            sr => \N__9514\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_57_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__10604\,
            in1 => \N__10100\,
            in2 => \_gnd_net_\,
            in3 => \N__8349\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9789\,
            ce => \N__9618\,
            sr => \N__9514\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_23_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__9183\,
            in1 => \N__10605\,
            in2 => \_gnd_net_\,
            in3 => \N__10101\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9789\,
            ce => \N__9618\,
            sr => \N__9514\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_27_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__10603\,
            in1 => \N__10099\,
            in2 => \_gnd_net_\,
            in3 => \N__6489\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9789\,
            ce => \N__9618\,
            sr => \N__9514\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_26_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__6495\,
            in1 => \N__10606\,
            in2 => \_gnd_net_\,
            in3 => \N__10102\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9789\,
            ce => \N__9618\,
            sr => \N__9514\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_60_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101010101111"
        )
    port map (
            in0 => \N__6483\,
            in1 => \_gnd_net_\,
            in2 => \N__10380\,
            in3 => \N__10682\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9785\,
            ce => \N__9614\,
            sr => \N__9518\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_61_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__10680\,
            in1 => \N__10289\,
            in2 => \_gnd_net_\,
            in3 => \N__6477\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9785\,
            ce => \N__9614\,
            sr => \N__9518\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_62_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__10681\,
            in1 => \N__10290\,
            in2 => \_gnd_net_\,
            in3 => \N__6471\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9785\,
            ce => \N__9614\,
            sr => \N__9518\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_30_LC_5_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__6990\,
            in1 => \N__10757\,
            in2 => \_gnd_net_\,
            in3 => \N__10319\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9781\,
            ce => \N__9610\,
            sr => \N__9522\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_31_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__6981\,
            in1 => \N__10758\,
            in2 => \_gnd_net_\,
            in3 => \N__10320\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9781\,
            ce => \N__9610\,
            sr => \N__9522\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_85_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__6677\,
            in1 => \N__6969\,
            in2 => \_gnd_net_\,
            in3 => \N__7707\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9816\,
            ce => \N__6578\,
            sr => \N__9493\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_84_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__6676\,
            in1 => \N__6975\,
            in2 => \_gnd_net_\,
            in3 => \N__7706\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9816\,
            ce => \N__6578\,
            sr => \N__9493\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_41_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__6821\,
            in1 => \N__6765\,
            in2 => \_gnd_net_\,
            in3 => \N__7695\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9811\,
            ce => \N__6579\,
            sr => \N__9497\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_87_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7693\,
            in1 => \N__6640\,
            in2 => \_gnd_net_\,
            in3 => \N__6585\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9811\,
            ce => \N__6579\,
            sr => \N__9497\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_40_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__6820\,
            in1 => \N__6774\,
            in2 => \_gnd_net_\,
            in3 => \N__7694\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9811\,
            ce => \N__6579\,
            sr => \N__9497\
        );

    \switch_clk_2MHz_inst.bit_sequence_stat_86_LC_6_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__7692\,
            in1 => \N__6639\,
            in2 => \_gnd_net_\,
            in3 => \N__6591\,
            lcout => \switch_clk_2MHz_inst.bit_sequence_statZ0Z_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9811\,
            ce => \N__6579\,
            sr => \N__9497\
        );

    \switch_clk_2MHz_inst.counter_din_RNO_0_2_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__7101\,
            in1 => \N__7048\,
            in2 => \N__7080\,
            in3 => \N__7155\,
            lcout => OPEN,
            ltout => \switch_clk_2MHz_inst.counter_din_3_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.counter_din_2_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__7400\,
            in1 => \N__7050\,
            in2 => \N__7116\,
            in3 => \N__7026\,
            lcout => \switch_clk_2MHz_inst.counter_dinZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9806\,
            ce => 'H',
            sr => \N__9500\
        );

    \switch_clk_2MHz_inst.counter_din_0_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__7102\,
            in1 => \N__7156\,
            in2 => \_gnd_net_\,
            in3 => \N__7399\,
            lcout => \switch_clk_2MHz_inst.counter_dinZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9806\,
            ce => 'H',
            sr => \N__9500\
        );

    \divisor_inst.clk_out_RNI3LEM_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8305\,
            in1 => \N__7288\,
            in2 => \_gnd_net_\,
            in3 => \N__8274\,
            lcout => \clk_out_RNI3LEM\,
            ltout => \clk_out_RNI3LEM_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.counter_din_1_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110000001100"
        )
    port map (
            in0 => \N__7103\,
            in1 => \N__7078\,
            in2 => \N__7113\,
            in3 => \N__7157\,
            lcout => \switch_clk_2MHz_inst.counter_dinZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9806\,
            ce => 'H',
            sr => \N__9500\
        );

    \switch_clk_2MHz_inst.current_state_RNO_5_0_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__7046\,
            in1 => \N__7070\,
            in2 => \N__7016\,
            in3 => \N__7099\,
            lcout => \switch_clk_2MHz_inst.G_31_0_o4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.counter_din_RNIBRN21_1_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__7100\,
            in1 => \_gnd_net_\,
            in2 => \N__7079\,
            in3 => \N__7047\,
            lcout => \switch_clk_2MHz_inst.N_92_0\,
            ltout => \switch_clk_2MHz_inst.N_92_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.counter_din_3_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110110000000"
        )
    port map (
            in0 => \N__7401\,
            in1 => \N__7158\,
            in2 => \N__7020\,
            in3 => \N__7015\,
            lcout => \switch_clk_2MHz_inst.counter_dinZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9806\,
            ce => 'H',
            sr => \N__9500\
        );

    \switch_clk_2MHz_inst.SEL_0_RNIC97Q_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__8275\,
            in1 => \N__7289\,
            in2 => \N__8315\,
            in3 => \N__7171\,
            lcout => \switch_clk_2MHz_inst.SEL_0_RNIC97QZ0\,
            ltout => \switch_clk_2MHz_inst.SEL_0_RNIC97QZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.SEL_0_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7317\,
            in2 => \N__6993\,
            in3 => \N__7153\,
            lcout => \switch_clk_2MHz_inst.aux_selection_2MHz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9802\,
            ce => 'H',
            sr => \N__9504\
        );

    \switch_clk_2MHz_inst.SEL_0_RNIC97Q_0_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100000000"
        )
    port map (
            in0 => \N__8277\,
            in1 => \N__7291\,
            in2 => \N__8316\,
            in3 => \N__7172\,
            lcout => \switch_clk_2MHz_inst.SEL_0_RNIC97QZ0Z_0\,
            ltout => \switch_clk_2MHz_inst.SEL_0_RNIC97QZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.SEL_0_RNILHTT1_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7152\,
            in2 => \N__7311\,
            in3 => \N__7308\,
            lcout => \N_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divisor_inst.clk_out_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__8278\,
            in1 => \N__8313\,
            in2 => \_gnd_net_\,
            in3 => \N__7292\,
            lcout => \clk_continuous_2MHz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9802\,
            ce => 'H',
            sr => \N__9504\
        );

    \switch_clk_2MHz_inst.current_state_fast_fast_RNITUE9_1_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7593\,
            in2 => \_gnd_net_\,
            in3 => \N__7214\,
            lcout => \switch_clk_2MHz_inst.N_91_li\,
            ltout => \switch_clk_2MHz_inst.N_91_li_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.current_state_fast_fast_RNI0KTV_1_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__8276\,
            in1 => \N__8312\,
            in2 => \N__7302\,
            in3 => \N__7290\,
            lcout => \switch_clk_2MHz_inst.current_state_fast_fast_RNI0KTVZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.current_state_fast_fast_1_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__7215\,
            in1 => \N__7594\,
            in2 => \N__7251\,
            in3 => \N__7402\,
            lcout => \switch_clk_2MHz_inst.current_state_fast_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9802\,
            ce => 'H',
            sr => \N__9504\
        );

    \mosi_output_obuf_RNO_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8155\,
            in1 => \N__9111\,
            in2 => \_gnd_net_\,
            in3 => \N__7203\,
            lcout => mosi_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.SEL_0_RNI98M31_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7173\,
            in2 => \N__7418\,
            in3 => \N__7154\,
            lcout => \switch_clk_2MHz_inst.SEL_0_RNI98MZ0Z31\,
            ltout => \switch_clk_2MHz_inst.SEL_0_RNI98MZ0Z31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.SEL_0_RNI4VEB3_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8458\,
            in2 => \N__7125\,
            in3 => \N__8168\,
            lcout => \N_381_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.SEL_0_er_RNIQKO61_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10264\,
            in1 => \N__8025\,
            in2 => \_gnd_net_\,
            in3 => \N__9076\,
            lcout => \N_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_2MHz_inst.flag_output_1_RNI12011_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__8154\,
            in1 => \N__7832\,
            in2 => \N__7490\,
            in3 => \N__7407\,
            lcout => \N_4_0\,
            ltout => \N_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_RNI7S8U1_15_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__8420\,
            in1 => \N__8408\,
            in2 => \N__8013\,
            in3 => \N__8841\,
            lcout => \delay_reg_RNI7S8U1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst.STATCNF_1_RNO_0_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__8010\,
            in1 => \N__8457\,
            in2 => \_gnd_net_\,
            in3 => \N__8001\,
            lcout => \config_register_latched_dec_inst.N_381_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_2_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8109\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9794\,
            ce => 'H',
            sr => \N__9510\
        );

    \divisor_inst_2.counter_2_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__8194\,
            in1 => \N__8235\,
            in2 => \_gnd_net_\,
            in3 => \N__8213\,
            lcout => \divisor_inst_2.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9794\,
            ce => 'H',
            sr => \N__9510\
        );

    \divisor_inst_2.counter_0_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8237\,
            lcout => \divisor_inst_2.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9794\,
            ce => 'H',
            sr => \N__9510\
        );

    \switch_clk_2MHz_inst.flag_output_1_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__8156\,
            in1 => \N__7831\,
            in2 => \N__7494\,
            in3 => \N__7411\,
            lcout => flag_signal,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9794\,
            ce => 'H',
            sr => \N__9510\
        );

    \divisor_inst_2.counter_1_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8193\,
            in2 => \_gnd_net_\,
            in3 => \N__8238\,
            lcout => \divisor_inst_2.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9794\,
            ce => 'H',
            sr => \N__9510\
        );

    \divisor_inst_2.clk_out_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__8236\,
            in1 => \N__8214\,
            in2 => \N__8199\,
            in3 => \N__8126\,
            lcout => \clk_continuous_1MHz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9794\,
            ce => 'H',
            sr => \N__9510\
        );

    \flag_output_ret_LC_6_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8175\,
            in1 => \N__8169\,
            in2 => \_gnd_net_\,
            in3 => \N__8459\,
            lcout => sel_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9794\,
            ce => 'H',
            sr => \N__9510\
        );

    \switch_clk_1MHz_inst.flag_input_reg_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8157\,
            lcout => \switch_clk_1MHz_inst.flag_input_regZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9790\,
            ce => 'H',
            sr => \N__9515\
        );

    \switch_clk_1MHz_inst.CLK_uC_LC_6_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011010010000"
        )
    port map (
            in0 => \N__10645\,
            in1 => \N__10218\,
            in2 => \N__8043\,
            in3 => \N__8127\,
            lcout => \switch_clk_1MHz_inst.CLK_uCZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9790\,
            ce => 'H',
            sr => \N__9515\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_1_LC_6_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8031\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9790\,
            ce => 'H',
            sr => \N__9515\
        );

    \switch_clk_1MHz_inst.counter_din_3_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110001000100"
        )
    port map (
            in0 => \N__9088\,
            in1 => \N__8060\,
            in2 => \N__8100\,
            in3 => \N__8088\,
            lcout => \switch_clk_1MHz_inst.counter_dinZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9790\,
            ce => 'H',
            sr => \N__9515\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_0_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8042\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9790\,
            ce => 'H',
            sr => \N__9515\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_64_LC_6_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__8337\,
            in1 => \N__10610\,
            in2 => \_gnd_net_\,
            in3 => \N__10260\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9786\,
            ce => \N__9615\,
            sr => \N__9519\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_55_LC_6_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__8496\,
            in1 => \N__10609\,
            in2 => \_gnd_net_\,
            in3 => \N__10259\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9786\,
            ce => \N__9615\,
            sr => \N__9519\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_56_LC_6_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10258\,
            in1 => \N__8355\,
            in2 => \_gnd_net_\,
            in3 => \N__10611\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9786\,
            ce => \N__9615\,
            sr => \N__9519\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_63_LC_6_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__8343\,
            in1 => \N__10891\,
            in2 => \_gnd_net_\,
            in3 => \N__10294\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9782\,
            ce => \N__9611\,
            sr => \N__9523\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_32_LC_6_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10890\,
            in1 => \N__8331\,
            in2 => \_gnd_net_\,
            in3 => \N__10318\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9778\,
            ce => \N__9608\,
            sr => \N__9527\
        );

    \CONSTANT_ONE_LUT4_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_6_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8244\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_reg_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9807\,
            ce => 'H',
            sr => \N__9501\
        );

    \divisor_inst.counter_1_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8279\,
            in2 => \_gnd_net_\,
            in3 => \N__8314\,
            lcout => divisor_inst_counter_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9803\,
            ce => 'H',
            sr => \N__9505\
        );

    \divisor_inst.counter_0_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8280\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => divisor_inst_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9803\,
            ce => 'H',
            sr => \N__9505\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_7_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8250\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9803\,
            ce => 'H',
            sr => \N__9505\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_5_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8484\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9803\,
            ce => 'H',
            sr => \N__9505\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_4_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8388\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9803\,
            ce => 'H',
            sr => \N__9505\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_8_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8478\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9803\,
            ce => 'H',
            sr => \N__9505\
        );

    \switch_clk_2MHz_inst.delay_inst.delay_reg_3_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8472\,
            lcout => \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9799\,
            ce => 'H',
            sr => \N__9508\
        );

    \flag_output_0_ret_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8409\,
            in1 => \N__8840\,
            in2 => \_gnd_net_\,
            in3 => \N__8460\,
            lcout => clk_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9799\,
            ce => 'H',
            sr => \N__9508\
        );

    \switch_clk_2MHz_inst.delay_inst.delay_reg_6_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8370\,
            lcout => \switch_clk_2MHz_inst_delay_inst_delay_reg_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9799\,
            ce => 'H',
            sr => \N__9508\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_3_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8397\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9799\,
            ce => 'H',
            sr => \N__9508\
        );

    \switch_clk_2MHz_inst.delay_inst.delay_reg_4_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8382\,
            lcout => \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9799\,
            ce => 'H',
            sr => \N__9508\
        );

    \switch_clk_2MHz_inst.delay_inst.delay_reg_5_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8376\,
            lcout => \switch_clk_2MHz_inst.delay_inst.delay_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9799\,
            ce => 'H',
            sr => \N__9508\
        );

    \config_register_latched_dec_inst.STATCNF_1_0_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__8707\,
            in1 => \N__8666\,
            in2 => \N__8804\,
            in3 => \N__8816\,
            lcout => \config_register_latched_dec_inst.STATCNF_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9795\,
            ce => \N__8364\,
            sr => \N__9511\
        );

    \config_register_latched_dec_inst.DYNSR_0_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8534\,
            in1 => \N__8704\,
            in2 => \_gnd_net_\,
            in3 => \N__8551\,
            lcout => \config_register_latched_dec_inst.DYNSRZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9791\,
            ce => \N__8517\,
            sr => \N__9516\
        );

    \config_register_latched_dec_inst.STATSR_0_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8703\,
            in1 => \N__8535\,
            in2 => \_gnd_net_\,
            in3 => \N__8665\,
            lcout => \config_register_latched_dec_inst.STATSRZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9791\,
            ce => \N__8517\,
            sr => \N__9516\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_12_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__8607\,
            in1 => \N__10646\,
            in2 => \_gnd_net_\,
            in3 => \N__10195\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9787\,
            ce => \N__9616\,
            sr => \N__9520\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_33_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10193\,
            in1 => \N__8505\,
            in2 => \_gnd_net_\,
            in3 => \N__10652\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9787\,
            ce => \N__9616\,
            sr => \N__9520\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_15_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__8625\,
            in1 => \N__10647\,
            in2 => \_gnd_net_\,
            in3 => \N__10196\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9787\,
            ce => \N__9616\,
            sr => \N__9520\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_54_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10194\,
            in1 => \N__8613\,
            in2 => \_gnd_net_\,
            in3 => \N__10653\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9787\,
            ce => \N__9616\,
            sr => \N__9520\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_52_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__8898\,
            in1 => \N__10648\,
            in2 => \_gnd_net_\,
            in3 => \N__10197\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9787\,
            ce => \N__9616\,
            sr => \N__9520\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_13_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10191\,
            in1 => \N__8490\,
            in2 => \_gnd_net_\,
            in3 => \N__10650\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9787\,
            ce => \N__9616\,
            sr => \N__9520\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_9_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__9225\,
            in1 => \N__10649\,
            in2 => \_gnd_net_\,
            in3 => \N__10198\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9787\,
            ce => \N__9616\,
            sr => \N__9520\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_14_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10192\,
            in1 => \N__8631\,
            in2 => \_gnd_net_\,
            in3 => \N__10651\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9787\,
            ce => \N__9616\,
            sr => \N__9520\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_53_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10769\,
            in1 => \N__8619\,
            in2 => \_gnd_net_\,
            in3 => \N__10263\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9783\,
            ce => \N__9612\,
            sr => \N__9524\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_11_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10261\,
            in1 => \N__8595\,
            in2 => \_gnd_net_\,
            in3 => \N__10770\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9783\,
            ce => \N__9612\,
            sr => \N__9524\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_10_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10768\,
            in1 => \N__8601\,
            in2 => \_gnd_net_\,
            in3 => \N__10262\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9783\,
            ce => \N__9612\,
            sr => \N__9524\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_13_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8562\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9796\,
            ce => 'H',
            sr => \N__9512\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_9_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8589\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9796\,
            ce => 'H',
            sr => \N__9512\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_11_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8574\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9796\,
            ce => 'H',
            sr => \N__9512\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_10_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8580\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9796\,
            ce => 'H',
            sr => \N__9512\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_12_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8568\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9796\,
            ce => 'H',
            sr => \N__9512\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_14_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8853\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_1MHz_inst.delay_inst.delay_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9792\,
            ce => 'H',
            sr => \N__9517\
        );

    \switch_clk_1MHz_inst.delay_inst.delay_reg_15_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8847\,
            lcout => \switch_clk_1MHz_inst_delay_inst_delay_reg_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9792\,
            ce => 'H',
            sr => \N__9517\
        );

    \config_register_latched_dec_inst.STATCNF_1_RNIRDN51_0_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__8820\,
            in1 => \N__8805\,
            in2 => \N__8726\,
            in3 => \N__8673\,
            lcout => \config_register_latched_dec_inst.STATCNF_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_81_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101010101111"
        )
    port map (
            in0 => \N__8991\,
            in1 => \_gnd_net_\,
            in2 => \N__10416\,
            in3 => \N__10916\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9784\,
            ce => \N__9613\,
            sr => \N__9525\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_50_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__10920\,
            in1 => \N__10389\,
            in2 => \_gnd_net_\,
            in3 => \N__8637\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9784\,
            ce => \N__9613\,
            sr => \N__9525\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_82_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__8649\,
            in1 => \_gnd_net_\,
            in2 => \N__10417\,
            in3 => \N__10917\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9784\,
            ce => \N__9613\,
            sr => \N__9525\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_87_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__10921\,
            in1 => \N__10390\,
            in2 => \_gnd_net_\,
            in3 => \N__8643\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9784\,
            ce => \N__9613\,
            sr => \N__9525\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_86_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__9021\,
            in1 => \_gnd_net_\,
            in2 => \N__10418\,
            in3 => \N__10918\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9784\,
            ce => \N__9613\,
            sr => \N__9525\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_49_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__10919\,
            in1 => \N__10388\,
            in2 => \_gnd_net_\,
            in3 => \N__8919\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9784\,
            ce => \N__9613\,
            sr => \N__9525\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_48_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__8934\,
            in1 => \_gnd_net_\,
            in2 => \N__10415\,
            in3 => \N__10915\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9784\,
            ce => \N__9613\,
            sr => \N__9525\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_16_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__8913\,
            in1 => \N__10878\,
            in2 => \_gnd_net_\,
            in3 => \N__10219\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9779\,
            ce => \N__9609\,
            sr => \N__9528\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_51_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__8904\,
            in1 => \N__10880\,
            in2 => \_gnd_net_\,
            in3 => \N__10221\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9779\,
            ce => \N__9609\,
            sr => \N__9528\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_35_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__8880\,
            in1 => \N__10879\,
            in2 => \_gnd_net_\,
            in3 => \N__10220\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9779\,
            ce => \N__9609\,
            sr => \N__9528\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_34_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__10876\,
            in1 => \N__10214\,
            in2 => \_gnd_net_\,
            in3 => \N__8889\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9779\,
            ce => \N__9609\,
            sr => \N__9528\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_66_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__8859\,
            in1 => \N__10881\,
            in2 => \_gnd_net_\,
            in3 => \N__10222\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9779\,
            ce => \N__9609\,
            sr => \N__9528\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_67_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__10877\,
            in1 => \N__10215\,
            in2 => \_gnd_net_\,
            in3 => \N__8874\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9779\,
            ce => \N__9609\,
            sr => \N__9528\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_42_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101010101111"
        )
    port map (
            in0 => \N__9198\,
            in1 => \_gnd_net_\,
            in2 => \N__10409\,
            in3 => \N__10909\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9776\,
            ce => \N__9606\,
            sr => \N__9530\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_74_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10912\,
            in1 => \N__9171\,
            in2 => \_gnd_net_\,
            in3 => \N__10351\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9776\,
            ce => \N__9606\,
            sr => \N__9530\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_65_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101010101111"
        )
    port map (
            in0 => \N__8868\,
            in1 => \_gnd_net_\,
            in2 => \N__10410\,
            in3 => \N__10910\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9776\,
            ce => \N__9606\,
            sr => \N__9530\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_76_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10914\,
            in1 => \N__8979\,
            in2 => \_gnd_net_\,
            in3 => \N__10353\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9776\,
            ce => \N__9606\,
            sr => \N__9530\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_75_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10913\,
            in1 => \N__8985\,
            in2 => \_gnd_net_\,
            in3 => \N__10352\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9776\,
            ce => \N__9606\,
            sr => \N__9530\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_68_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101010101111"
        )
    port map (
            in0 => \N__8973\,
            in1 => \_gnd_net_\,
            in2 => \N__10411\,
            in3 => \N__10911\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9776\,
            ce => \N__9606\,
            sr => \N__9530\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_46_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100100001001000"
        )
    port map (
            in0 => \N__10374\,
            in1 => \N__8946\,
            in2 => \N__10966\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9774\,
            ce => \N__9604\,
            sr => \N__9533\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_43_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__8964\,
            in1 => \N__10922\,
            in2 => \_gnd_net_\,
            in3 => \N__10376\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9774\,
            ce => \N__9604\,
            sr => \N__9533\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_44_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110110111101101"
        )
    port map (
            in0 => \N__10373\,
            in1 => \N__8958\,
            in2 => \N__10965\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9774\,
            ce => \N__9604\,
            sr => \N__9533\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_45_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__8952\,
            in1 => \N__10923\,
            in2 => \_gnd_net_\,
            in3 => \N__10377\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9774\,
            ce => \N__9604\,
            sr => \N__9533\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_47_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__8940\,
            in1 => \N__10924\,
            in2 => \_gnd_net_\,
            in3 => \N__10378\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9774\,
            ce => \N__9604\,
            sr => \N__9533\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_69_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100100001001000"
        )
    port map (
            in0 => \N__10375\,
            in1 => \N__8925\,
            in2 => \N__10967\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9774\,
            ce => \N__9604\,
            sr => \N__9533\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_70_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__9147\,
            in1 => \N__10934\,
            in2 => \_gnd_net_\,
            in3 => \N__10386\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9771\,
            ce => \N__9601\,
            sr => \N__9536\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_71_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__9141\,
            in1 => \N__10935\,
            in2 => \_gnd_net_\,
            in3 => \N__10387\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9771\,
            ce => \N__9601\,
            sr => \N__9536\
        );

    \switch_clk_1MHz_inst.MOSI_er_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__9135\,
            in1 => \N__10941\,
            in2 => \N__9123\,
            in3 => \N__10372\,
            lcout => \mosi_1MHz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9780\,
            ce => \N__9102\,
            sr => \N__9521\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_85_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__10939\,
            in1 => \N__10404\,
            in2 => \_gnd_net_\,
            in3 => \N__9003\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9777\,
            ce => \N__9607\,
            sr => \N__9526\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_83_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__9015\,
            in1 => \_gnd_net_\,
            in2 => \N__10419\,
            in3 => \N__10940\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9777\,
            ce => \N__9607\,
            sr => \N__9526\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_84_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__10938\,
            in1 => \N__10403\,
            in2 => \_gnd_net_\,
            in3 => \N__9009\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9777\,
            ce => \N__9607\,
            sr => \N__9526\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_17_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__8997\,
            in1 => \N__10882\,
            in2 => \_gnd_net_\,
            in3 => \N__10203\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9775\,
            ce => \N__9605\,
            sr => \N__9529\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_40_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10199\,
            in1 => \N__9240\,
            in2 => \_gnd_net_\,
            in3 => \N__10886\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9775\,
            ce => \N__9605\,
            sr => \N__9529\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_80_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__9291\,
            in1 => \N__10885\,
            in2 => \_gnd_net_\,
            in3 => \N__10206\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9775\,
            ce => \N__9605\,
            sr => \N__9529\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_8_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10202\,
            in1 => \N__9216\,
            in2 => \_gnd_net_\,
            in3 => \N__10889\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9775\,
            ce => \N__9605\,
            sr => \N__9529\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_7_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__9210\,
            in1 => \N__10884\,
            in2 => \_gnd_net_\,
            in3 => \N__10205\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9775\,
            ce => \N__9605\,
            sr => \N__9529\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_6_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10201\,
            in1 => \N__9279\,
            in2 => \_gnd_net_\,
            in3 => \N__10888\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9775\,
            ce => \N__9605\,
            sr => \N__9529\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_21_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__9153\,
            in1 => \N__10883\,
            in2 => \_gnd_net_\,
            in3 => \N__10204\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9775\,
            ce => \N__9605\,
            sr => \N__9529\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_41_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10200\,
            in1 => \N__9204\,
            in2 => \_gnd_net_\,
            in3 => \N__10887\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9775\,
            ce => \N__9605\,
            sr => \N__9529\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_22_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10937\,
            in1 => \N__9192\,
            in2 => \_gnd_net_\,
            in3 => \N__10363\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9772\,
            ce => \N__9602\,
            sr => \N__9531\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_73_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__9159\,
            in1 => \N__10905\,
            in2 => \_gnd_net_\,
            in3 => \N__10379\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9769\,
            ce => \N__9599\,
            sr => \N__9534\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_72_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10385\,
            in1 => \N__9165\,
            in2 => \_gnd_net_\,
            in3 => \N__10936\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9766\,
            ce => \N__9596\,
            sr => \N__9537\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_20_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100100001001000"
        )
    port map (
            in0 => \N__10207\,
            in1 => \N__9267\,
            in2 => \N__10968\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9773\,
            ce => \N__9603\,
            sr => \N__9532\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_18_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__9303\,
            in1 => \N__10948\,
            in2 => \_gnd_net_\,
            in3 => \N__10211\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9773\,
            ce => \N__9603\,
            sr => \N__9532\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_4_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100100001001000"
        )
    port map (
            in0 => \N__10208\,
            in1 => \N__9231\,
            in2 => \N__10969\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9773\,
            ce => \N__9603\,
            sr => \N__9532\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_78_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__9249\,
            in1 => \N__10950\,
            in2 => \_gnd_net_\,
            in3 => \N__10213\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9773\,
            ce => \N__9603\,
            sr => \N__9532\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_79_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100100001001000"
        )
    port map (
            in0 => \N__10210\,
            in1 => \N__9297\,
            in2 => \N__10971\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9773\,
            ce => \N__9603\,
            sr => \N__9532\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_5_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110110111101101"
        )
    port map (
            in0 => \N__10209\,
            in1 => \N__9285\,
            in2 => \N__10970\,
            in3 => \_gnd_net_\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9773\,
            ce => \N__9603\,
            sr => \N__9532\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_19_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__9273\,
            in1 => \N__10949\,
            in2 => \_gnd_net_\,
            in3 => \N__10212\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9773\,
            ce => \N__9603\,
            sr => \N__9532\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_77_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__9261\,
            in1 => \N__10906\,
            in2 => \_gnd_net_\,
            in3 => \N__10414\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9767\,
            ce => \N__9597\,
            sr => \N__9538\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_39_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__10945\,
            in1 => \N__10217\,
            in2 => \_gnd_net_\,
            in3 => \N__11013\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9770\,
            ce => \N__9600\,
            sr => \N__9535\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_3_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__11007\,
            in1 => \N__10947\,
            in2 => \_gnd_net_\,
            in3 => \N__10224\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9770\,
            ce => \N__9600\,
            sr => \N__9535\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_38_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__10944\,
            in1 => \N__10216\,
            in2 => \_gnd_net_\,
            in3 => \N__10986\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9770\,
            ce => \N__9600\,
            sr => \N__9535\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_2_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__10995\,
            in1 => \N__10946\,
            in2 => \_gnd_net_\,
            in3 => \N__10223\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9770\,
            ce => \N__9600\,
            sr => \N__9535\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_0_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10907\,
            in2 => \_gnd_net_\,
            in3 => \N__10413\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9765\,
            ce => \N__9595\,
            sr => \N__9540\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_1_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__10412\,
            in1 => \N__11001\,
            in2 => \_gnd_net_\,
            in3 => \N__10908\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9765\,
            ce => \N__9595\,
            sr => \N__9540\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_37_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__9840\,
            in1 => \N__10943\,
            in2 => \_gnd_net_\,
            in3 => \N__10226\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9768\,
            ce => \N__9598\,
            sr => \N__9539\
        );

    \switch_clk_1MHz_inst.bit_sequence_stat_36_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__10980\,
            in1 => \N__10942\,
            in2 => \_gnd_net_\,
            in3 => \N__10225\,
            lcout => \switch_clk_1MHz_inst.bit_sequence_statZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9768\,
            ce => \N__9598\,
            sr => \N__9539\
        );

    \config_register_latched_dec_inst.STATCNF_1_RNIRDN51_0_0_LC_32_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9324\,
            lcout => \STATCNF_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
